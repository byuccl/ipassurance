module graphiti
   (clk,
    clk15M,
    reset,
    \output ,
    in_r,
    in_g,
    in_b,
    framereset,
    en_bild,
    readmem);
  input clk;
  input clk15M;
  input reset;
  output [15:0]\output ;
  input [4:0]in_r;
  input [4:0]in_g;
  input [4:0]in_b;
  output framereset;
  output en_bild;
  output readmem;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]A;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [22:1]C;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [22:1]C__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire GND_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild12_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_bild1_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_burst0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_burst1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/en_burst10_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\I_0/hlctr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr2_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/hlctr_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_austastung ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_austastung1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_austastung2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_sync_last ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_vertbr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_vertbr1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_vertbr131_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_vertbr2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_vertbr_last ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_verteq1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_en_verteq2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_framereset ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase433_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_phase4_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_readmem1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_readmem15_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_readmem2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_readmem26_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]\I_0/i_sync_c ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c210_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c211_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c212_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c213_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c215_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c216_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c218_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c219_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c221_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c223_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c224_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c226_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c227_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c229_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c28_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/i_sync_c2_inferred__9_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/p_1_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\I_0/pixctr ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr1_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__6_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__6_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__6_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry__6_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr2_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_0/pixctr_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/abschnittu_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/adr_reg_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:1]\I_1/ctr90_48_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:1]\I_1/ctr_48_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_1/data_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_10 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_11 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_12 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_13 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_14 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_16 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_18 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_19 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_21 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_22 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_23 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_24 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_25 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_26 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_27 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_28 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_29 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_30 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_31 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_8 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/adr_reg_n_9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_2/data[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_CARRY4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_CARRY4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_CARRY4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/minusOp_inferred__0_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp__0_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/multOp_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/out_y_reg_c_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_3/plusOp__0_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\I_4/multOp__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp__39_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/multOp_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/output_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__2_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp__3_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__3_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__5_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__6_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7__62_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_inferred__7_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_4/plusOp_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\I_5/multOp__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp__39_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/multOp_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/output_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__0_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__1_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__2_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_100 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_101 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_102 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_103 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_104 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_105 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_58 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_59 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_60 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_61 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_62 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_63 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_64 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_65 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_66 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_67 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_68 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_69 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_70 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_71 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_72 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_73 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_74 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_77 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_78 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_79 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_80 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_81 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_82 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_84 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_85 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_86 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_87 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_88 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_89 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_90 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_91 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_93 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_94 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_96 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_97 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_98 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp__3_n_99 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__3_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__5_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__6_carry_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry__4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7__62_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry__4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_inferred__7_carry_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_106 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_108 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_109 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_110 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_111 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_112 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_113 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_115 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_116 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_117 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_118 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_119 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_120 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_121 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_123 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_125 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_126 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_127 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_129 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_130 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_131 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_132 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_133 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_134 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_135 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_136 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_137 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_138 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_139 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_140 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_141 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_142 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_143 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_144 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_145 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_146 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_147 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_148 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_149 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_150 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_151 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/plusOp_n_153 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[0][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[10][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[11][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[12][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[13][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[14][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[1][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[2][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[3][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[4][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[5][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[6][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[7][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[8][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_5/sr_reg_n_0_[9][9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/output_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][10]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][1]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][2]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][3]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][4]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][5]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][6]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][7]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][8]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[5][9]_srl7_I_6_sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][0]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][10]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][1]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][2]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][3]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][4]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][5]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][6]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][7]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][8]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg[6][9]_I_6_sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_c_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \I_6/sr_reg_gate_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]L;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]R;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire VCC_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire abschnittu;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \abschnittu[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \abschnittu[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \abschnittu[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \abschnittu[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]abschnittu_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_100_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_101_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_102_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_102_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_102_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_102_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_106_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_107_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_107_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_107_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_107_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_111_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_112_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_112_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_112_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_112_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_116_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_117_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_117_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_117_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_117_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_121_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_122_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_122_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_122_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_122_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_124_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_125_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_126_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_127_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_127_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_127_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_127_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_129_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_130_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_131_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_132_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_132_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_132_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_132_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_134_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_137_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_137_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_137_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_137_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_139_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_142_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_142_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_142_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_142_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_143_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_144_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_145_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_146_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_147_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_147_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_147_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_147_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_148_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_149_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_150_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_151_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_154_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_157_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_15_n_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_16_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_16_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_16_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_17_n_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_18_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_18_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_18_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_27_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_27_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_27_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_32_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_32_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_32_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_37_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_37_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_37_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_42_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_42_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_42_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_47_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_47_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_47_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_52_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_52_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_52_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_57_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_57_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_57_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_62_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_62_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_62_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_67_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_67_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_67_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_68_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_69_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_70_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_72_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_72_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_72_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_72_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_77_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_77_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_77_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_77_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_82_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_82_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_82_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_82_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_84_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_86_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_87_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_87_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_87_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_87_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_89_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_91_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_92_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_92_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_92_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_92_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_95_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_96_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_97_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_97_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_97_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire adr_reg_i_97_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire austastung_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clear;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk15M;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ctr90_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[37]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[41]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[45]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[45]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[45]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[49]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[53]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]ctr90_48_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[13]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[13]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[13]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[13]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[17]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[1]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[21]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[25]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[29]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[33]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[37]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[41]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[45]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[49]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[53]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[57]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[5]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[61]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[61]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[61]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[61]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr90_48_reg[9]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ctr_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[37]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[41]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[45]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[45]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[45]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[49]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[53]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]ctr_48_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[13]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[13]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[13]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[13]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[17]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[1]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[21]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[25]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[29]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[33]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[37]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[41]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[45]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[49]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[53]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[57]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[5]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[61]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[61]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[61]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[61]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \ctr_48_reg[9]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:1]data0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]data_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[12]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[15]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[4]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2__0_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \data_reg[8]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry__2_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild1_inferred__0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_10_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_10_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_10_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_15_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_15_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_15_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_3_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_3_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_3_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_bild_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_10_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_10_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_10_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_19_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_19_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_19_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_24_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_24_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_24_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_2_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_2_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_2_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_33_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_33_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_33_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_38_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_38_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_38_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_3_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_3_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_3_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire en_burst_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire framereset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire framereset_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0__0__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b9__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire g0_b9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire hlctr1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_12_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_12_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_12_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_18_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_18_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_18_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_23_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_23_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_23_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_28_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_28_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_28_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_34_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_34_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_34_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_5_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_5_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_5_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_6_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_6_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_austastung_reg_i_6_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_14_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_14_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_14_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_2_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_2_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_2_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_3_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_3_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_3_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_9_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_9_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_sync_last_reg_i_9_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_66_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_68_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_69_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_70_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_71_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_72_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_73_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_74_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_75_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_76_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_77_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_78_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_79_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_80_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_81_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_82_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_83_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_84_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_85_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_86_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_11_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_11_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_11_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_17_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_17_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_17_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_26_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_26_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_26_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_2_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_2_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_2_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_31_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_31_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_31_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_36_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_36_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_36_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_3_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_3_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_3_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_45_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_45_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_45_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_51_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_51_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_51_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_57_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_57_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_57_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_5_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_5_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_en_vertbr_last_reg_i_5_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry__2_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase4_inferred__0_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_phase_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_100_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_101_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_102_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_103_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_104_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_105_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_106_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_107_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_108_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_109_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_110_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_111_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_112_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_113_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_114_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_115_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_116_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_117_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_118_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_119_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_120_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_121_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_122_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_123_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_124_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_62_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_66_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_68_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_69_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_70_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_71_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_72_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_74_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_75_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_76_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_77_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_78_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_80_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_81_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_82_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_83_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_84_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_85_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_86_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_87_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_89_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_90_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_91_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_92_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_93_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_94_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_95_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_96_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_97_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_98_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_99_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_15_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_15_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_15_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_21_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_21_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_21_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_2_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_2_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_2_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_30_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_30_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_30_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_36_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_36_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_36_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_3_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_3_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_3_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_45_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_45_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_45_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_50_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_50_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_50_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_59_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_59_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_59_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_5_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_5_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_5_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_64_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_64_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_64_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_6_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_6_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_6_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_73_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_73_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_73_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_73_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_79_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_79_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_79_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_79_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_88_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_88_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_88_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_readmem_reg_i_88_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry__2_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_sync_c2_inferred__9_carry_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_119_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_121_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_122_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_123_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_124_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_125_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_127_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_128_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_129_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_130_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_131_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_132_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_133_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_134_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_136_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_137_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_138_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_139_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_145_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_146_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_147_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_148_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_150_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_151_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_152_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_153_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_155_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_156_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_157_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_158_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_159_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_160_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_161_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_162_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_164_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_165_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_166_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_167_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_168_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_169_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_170_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_171_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_173_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_174_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_175_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_176_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_177_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_178_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_179_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_180_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_182_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_183_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_184_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_185_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_187_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_188_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_189_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_190_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_192_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_193_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_194_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_195_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_196_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_197_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_198_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_199_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_201_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_202_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_203_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_204_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_206_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_207_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_208_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_209_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_210_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_211_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_212_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_213_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_215_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_216_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_217_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_218_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_220_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_221_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_222_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_223_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_224_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_225_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_226_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_227_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_229_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_230_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_231_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_232_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_234_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_235_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_236_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_237_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_238_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_239_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_240_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_241_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_243_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_244_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_245_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_246_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_248_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_249_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_250_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_251_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_252_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_253_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_254_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_255_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_257_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_258_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_259_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_260_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_261_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_263_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_264_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_265_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_266_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_267_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_268_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_269_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_270_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_272_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_273_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_274_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_275_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_276_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_277_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_278_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_279_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_281_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_282_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_283_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_284_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_285_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_286_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_287_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_288_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_290_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_291_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_292_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_293_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_294_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_296_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_297_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_298_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_299_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_300_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_302_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_303_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_304_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_305_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_306_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_307_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_308_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_309_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_311_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_312_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_313_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_314_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_315_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_317_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_318_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_319_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_320_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_321_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_322_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_323_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_324_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_326_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_327_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_328_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_329_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_330_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_332_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_333_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_334_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_335_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_336_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_337_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_338_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_339_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_341_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_342_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_343_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_344_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_346_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_347_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_348_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_349_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_350_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_351_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_352_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_353_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_354_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_355_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_356_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_357_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_358_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_359_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_360_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_361_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_362_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_363_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_364_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_365_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_366_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_367_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_368_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_369_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_370_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_371_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_372_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_373_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_374_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_375_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_376_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_377_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_378_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_379_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_380_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_381_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_382_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_383_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_384_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_385_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_386_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_387_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_388_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_389_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_390_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_391_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_392_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_393_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_394_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_395_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_396_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_397_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_398_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_399_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_400_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_401_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_402_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_403_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_404_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_405_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_406_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_407_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_408_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_409_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_410_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_411_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_412_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_413_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_414_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_415_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_416_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_417_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_418_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_419_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_420_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_421_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_422_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_423_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_424_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_425_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_426_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_427_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_428_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_429_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_430_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_431_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_432_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_433_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_434_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_435_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_436_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_437_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_438_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_439_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_440_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_441_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_442_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_443_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_444_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_445_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_446_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_447_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_448_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_449_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_450_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_451_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_452_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_453_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_454_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_455_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_456_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_457_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c[1]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]i_sync_c_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_111_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_111_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_111_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_120_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_120_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_120_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_120_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_126_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_126_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_126_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_126_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_135_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_135_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_135_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_135_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_140_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_140_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_140_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_140_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_149_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_149_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_149_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_149_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_154_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_154_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_154_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_154_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_163_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_163_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_163_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_163_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_16_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_172_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_172_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_172_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_172_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_181_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_181_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_181_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_181_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_186_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_186_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_186_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_186_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_191_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_191_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_191_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_191_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_200_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_200_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_200_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_200_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_205_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_205_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_205_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_205_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_214_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_214_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_214_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_214_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_219_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_219_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_219_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_219_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_21_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_21_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_21_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_228_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_228_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_228_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_228_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_233_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_233_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_233_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_233_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_242_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_242_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_242_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_242_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_247_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_247_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_247_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_247_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_256_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_256_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_256_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_256_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_262_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_262_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_262_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_262_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_271_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_271_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_271_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_271_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_27_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_27_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_27_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_280_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_280_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_280_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_280_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_289_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_289_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_289_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_289_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_295_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_295_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_295_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_295_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_301_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_301_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_301_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_301_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_310_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_310_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_310_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_310_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_316_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_316_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_316_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_316_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_325_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_325_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_325_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_325_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_331_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_331_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_331_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_331_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_340_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_340_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_340_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_340_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_345_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_345_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_345_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_345_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_36_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_36_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_36_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_42_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_42_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_42_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_51_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_51_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_51_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_60_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_60_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_60_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_69_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_69_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_69_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_75_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_75_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_75_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_81_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_81_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_81_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_90_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_90_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_90_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_96_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_96_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_96_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_sync_c_reg[1]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]in_b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]in_g;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]in_r;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\input ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire lopt;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire minusOp_inferred__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_100;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_101;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_102;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_103;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_104;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_105;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_64;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_65;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_67;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_68;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_69;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_70;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_71;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_72;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_73;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_74;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_75;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_76;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_77;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_78;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_79;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_80;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_81;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_82;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_83;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_84;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_85;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_86;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_87;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_88;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_89;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_90;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_91;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_92;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_93;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_94;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_95;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_96;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_97;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_98;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modu_reg_n_99;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_100;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_101;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_102;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_103;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_104;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_105;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_64;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_65;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_67;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_68;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_69;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_70;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_71;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_72;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_73;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_74;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_75;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_76;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_77;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_78;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_79;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_96;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_97;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_98;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modus_reg_n_99;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_16_n_4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_17_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_17_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_17_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_18_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_18_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_18_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_19_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_19_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_19_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_100;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_101;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_102;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_103;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_104;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_105;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_64;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_65;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_67;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_68;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_69;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_70;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_71;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_72;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_73;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_74;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_75;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_76;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_77;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_78;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_91;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_92;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_93;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_94;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_95;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_96;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_97;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_98;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modv_reg_n_99;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_100;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_101;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_102;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_103;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_104;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_105;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_64;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_65;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_67;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_68;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_69;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_70;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_71;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_72;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_73;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_74;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_75;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_76;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_77;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_78;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_79;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_96;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_97;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_98;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modvs_reg_n_99;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_100;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_101;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_102;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_103;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_104;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_105;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_58;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_59;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_60;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_61;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_62;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_63;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_64;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_65;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_67;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_68;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_69;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_70;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_71;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_72;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_73;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_74;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_75;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_76;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_77;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_78;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_79;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_80;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_81;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_82;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_83;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_84;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_85;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_86;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_87;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_88;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_89;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_90;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_91;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_92;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_93;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_94;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_95;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_96;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_97;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_98;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire modys_reg_n_99;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]multOp0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_8__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__1_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_6__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_7__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp__39_carry_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire multOp_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]\output ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]output_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[0]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[12]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[15]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[4]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \output_reg[8]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]p_1_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_2_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]p_2_in__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_3_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [7:0]p_3_in__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire phase;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire pixctr1_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]plusOp0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [10:0]plusOp18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__0_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp__0_carry_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__3_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__5_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__6_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__2_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__3_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry__4_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7__62_carry_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__0_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__1_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_5__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__2_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_4__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__3_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__4_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__4_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__4_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry__4_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_2__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_3__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire plusOp_inferred__7_carry_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]pre_yuv_v;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:0]prevideo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:1]psin0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire readmem;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sr;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \sr[2][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sr_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\sr_reg[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_12_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_12_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_12_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_18_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_18_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_18_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_23_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_23_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_23_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_28_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_28_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_28_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_33_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_33_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_33_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_4_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_4_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_4_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_5_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_5_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_5_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_6_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_6_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire sync_reg_i_6_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tmr_austastung;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire tmr_en_burst;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_1
       (.G(GND_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/austastung_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(austastung_i_1_n_0),
        .Q(tmr_austastung));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/en_bild1_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/en_bild1_inferred__0_carry_n_0 ,\I_0/en_bild1_inferred__0_carry_n_1 ,\I_0/en_bild1_inferred__0_carry_n_2 ,\I_0/en_bild1_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({en_bild1_inferred__0_carry_i_1_n_0,en_bild1_inferred__0_carry_i_2_n_0,\<const0>__0__0 ,en_bild1_inferred__0_carry_i_3_n_0}),
        .S({en_bild1_inferred__0_carry_i_4_n_0,en_bild1_inferred__0_carry_i_5_n_0,en_bild1_inferred__0_carry_i_6_n_0,en_bild1_inferred__0_carry_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/en_bild1_inferred__0_carry__0 
       (.CI(\I_0/en_bild1_inferred__0_carry_n_0 ),
        .CO({\I_0/en_bild1_inferred__0_carry__0_n_0 ,\I_0/en_bild1_inferred__0_carry__0_n_1 ,\I_0/en_bild1_inferred__0_carry__0_n_2 ,\I_0/en_bild1_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_bild1_inferred__0_carry__0_i_1_n_0,en_bild1_inferred__0_carry__0_i_2_n_0,en_bild1_inferred__0_carry__0_i_3_n_0,en_bild1_inferred__0_carry__0_i_4_n_0}),
        .S({en_bild1_inferred__0_carry__0_i_5_n_0,en_bild1_inferred__0_carry__0_i_6_n_0,en_bild1_inferred__0_carry__0_i_7_n_0,en_bild1_inferred__0_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/en_bild1_inferred__0_carry__1 
       (.CI(\I_0/en_bild1_inferred__0_carry__0_n_0 ),
        .CO({\I_0/en_bild1_inferred__0_carry__1_n_0 ,\I_0/en_bild1_inferred__0_carry__1_n_1 ,\I_0/en_bild1_inferred__0_carry__1_n_2 ,\I_0/en_bild1_inferred__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_bild1_inferred__0_carry__1_i_1_n_0,en_bild1_inferred__0_carry__1_i_2_n_0,en_bild1_inferred__0_carry__1_i_3_n_0,en_bild1_inferred__0_carry__1_i_4_n_0}),
        .S({en_bild1_inferred__0_carry__1_i_5_n_0,en_bild1_inferred__0_carry__1_i_6_n_0,en_bild1_inferred__0_carry__1_i_7_n_0,en_bild1_inferred__0_carry__1_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/en_bild1_inferred__0_carry__2 
       (.CI(\I_0/en_bild1_inferred__0_carry__1_n_0 ),
        .CO({\I_0/en_bild12_in ,\I_0/en_bild1_inferred__0_carry__2_n_1 ,\I_0/en_bild1_inferred__0_carry__2_n_2 ,\I_0/en_bild1_inferred__0_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_bild1_inferred__0_carry__2_i_1_n_0,en_bild1_inferred__0_carry__2_i_2_n_0,en_bild1_inferred__0_carry__2_i_3_n_0,en_bild1_inferred__0_carry__2_i_4_n_0}),
        .S({en_bild1_inferred__0_carry__2_i_5_n_0,en_bild1_inferred__0_carry__2_i_6_n_0,en_bild1_inferred__0_carry__2_i_7_n_0,en_bild1_inferred__0_carry__2_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/en_bild_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_0/en_bild0 ),
        .Q(en_bild));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/en_burst_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_0/en_burst0 ),
        .Q(tmr_en_burst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_0/framereset_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(framereset_i_1_n_0),
        .PRE(clear),
        .Q(framereset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/hlctr1_carry_n_0 ,\I_0/hlctr1_carry_n_1 ,\I_0/hlctr1_carry_n_2 ,\I_0/hlctr1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({hlctr1_carry_i_1_n_0,hlctr1_carry_i_2_n_0,hlctr1_carry_i_3_n_0,hlctr1_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr1_carry__0 
       (.CI(\I_0/hlctr1_carry_n_0 ),
        .CO({\I_0/hlctr1_carry__0_n_0 ,\I_0/hlctr1_carry__0_n_1 ,\I_0/hlctr1_carry__0_n_2 ,\I_0/hlctr1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({hlctr1_carry__0_i_1_n_0,hlctr1_carry__0_i_2_n_0,hlctr1_carry__0_i_3_n_0,hlctr1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr1_carry__1 
       (.CI(\I_0/hlctr1_carry__0_n_0 ),
        .CO({\I_0/hlctr1_carry__1_n_0 ,\I_0/hlctr1_carry__1_n_1 ,\I_0/hlctr1_carry__1_n_2 ,\I_0/hlctr1_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,hlctr1_carry__1_i_1_n_0,hlctr1_carry__1_i_2_n_0,hlctr1_carry__1_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/hlctr2_carry_n_0 ,\I_0/hlctr2_carry_n_1 ,\I_0/hlctr2_carry_n_2 ,\I_0/hlctr2_carry_n_3 }),
        .CYINIT(\I_0/hlctr_reg_n_0_ ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry_n_4 ,\I_0/hlctr2_carry_n_5 ,\I_0/hlctr2_carry_n_6 ,\I_0/hlctr2_carry_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[4] ,\I_0/hlctr_reg_n_0_[3] ,\I_0/hlctr_reg_n_0_[2] ,\I_0/hlctr_reg_n_0_[1] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__0 
       (.CI(\I_0/hlctr2_carry_n_0 ),
        .CO({\I_0/hlctr2_carry__0_n_0 ,\I_0/hlctr2_carry__0_n_1 ,\I_0/hlctr2_carry__0_n_2 ,\I_0/hlctr2_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__0_n_4 ,\I_0/hlctr2_carry__0_n_5 ,\I_0/hlctr2_carry__0_n_6 ,\I_0/hlctr2_carry__0_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[8] ,\I_0/hlctr_reg_n_0_[7] ,\I_0/hlctr_reg_n_0_[6] ,\I_0/hlctr_reg_n_0_[5] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__1 
       (.CI(\I_0/hlctr2_carry__0_n_0 ),
        .CO({\I_0/hlctr2_carry__1_n_0 ,\I_0/hlctr2_carry__1_n_1 ,\I_0/hlctr2_carry__1_n_2 ,\I_0/hlctr2_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__1_n_4 ,\I_0/hlctr2_carry__1_n_5 ,\I_0/hlctr2_carry__1_n_6 ,\I_0/hlctr2_carry__1_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[12] ,\I_0/hlctr_reg_n_0_[11] ,\I_0/hlctr_reg_n_0_[10] ,\I_0/hlctr_reg_n_0_[9] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__2 
       (.CI(\I_0/hlctr2_carry__1_n_0 ),
        .CO({\I_0/hlctr2_carry__2_n_0 ,\I_0/hlctr2_carry__2_n_1 ,\I_0/hlctr2_carry__2_n_2 ,\I_0/hlctr2_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__2_n_4 ,\I_0/hlctr2_carry__2_n_5 ,\I_0/hlctr2_carry__2_n_6 ,\I_0/hlctr2_carry__2_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[16] ,\I_0/hlctr_reg_n_0_[15] ,\I_0/hlctr_reg_n_0_[14] ,\I_0/hlctr_reg_n_0_[13] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__3 
       (.CI(\I_0/hlctr2_carry__2_n_0 ),
        .CO({\I_0/hlctr2_carry__3_n_0 ,\I_0/hlctr2_carry__3_n_1 ,\I_0/hlctr2_carry__3_n_2 ,\I_0/hlctr2_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__3_n_4 ,\I_0/hlctr2_carry__3_n_5 ,\I_0/hlctr2_carry__3_n_6 ,\I_0/hlctr2_carry__3_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[20] ,\I_0/hlctr_reg_n_0_[19] ,\I_0/hlctr_reg_n_0_[18] ,\I_0/hlctr_reg_n_0_[17] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__4 
       (.CI(\I_0/hlctr2_carry__3_n_0 ),
        .CO({\I_0/hlctr2_carry__4_n_0 ,\I_0/hlctr2_carry__4_n_1 ,\I_0/hlctr2_carry__4_n_2 ,\I_0/hlctr2_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__4_n_4 ,\I_0/hlctr2_carry__4_n_5 ,\I_0/hlctr2_carry__4_n_6 ,\I_0/hlctr2_carry__4_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[24] ,\I_0/hlctr_reg_n_0_[23] ,\I_0/hlctr_reg_n_0_[22] ,\I_0/hlctr_reg_n_0_[21] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__5 
       (.CI(\I_0/hlctr2_carry__4_n_0 ),
        .CO({\I_0/hlctr2_carry__5_n_0 ,\I_0/hlctr2_carry__5_n_1 ,\I_0/hlctr2_carry__5_n_2 ,\I_0/hlctr2_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__5_n_4 ,\I_0/hlctr2_carry__5_n_5 ,\I_0/hlctr2_carry__5_n_6 ,\I_0/hlctr2_carry__5_n_7 }),
        .S({\I_0/hlctr_reg_n_0_[28] ,\I_0/hlctr_reg_n_0_[27] ,\I_0/hlctr_reg_n_0_[26] ,\I_0/hlctr_reg_n_0_[25] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/hlctr2_carry__6 
       (.CI(\I_0/hlctr2_carry__5_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/hlctr2_carry__6_n_4 ,\I_0/hlctr2_carry__6_n_5 ,\I_0/hlctr2_carry__6_n_6 ,\I_0/hlctr2_carry__6_n_7 }),
        .S({\<const0>__0__0 ,\I_0/hlctr_reg_n_0_[31] ,\I_0/hlctr_reg_n_0_[30] ,\I_0/hlctr_reg_n_0_[29] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[0] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [0]),
        .Q(\I_0/hlctr_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[10] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [10]),
        .Q(\I_0/hlctr_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[11] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [11]),
        .Q(\I_0/hlctr_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[12] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [12]),
        .Q(\I_0/hlctr_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[13] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [13]),
        .Q(\I_0/hlctr_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[14] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [14]),
        .Q(\I_0/hlctr_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[15] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [15]),
        .Q(\I_0/hlctr_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[16] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [16]),
        .Q(\I_0/hlctr_reg_n_0_[16] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[17] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [17]),
        .Q(\I_0/hlctr_reg_n_0_[17] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[18] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [18]),
        .Q(\I_0/hlctr_reg_n_0_[18] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[19] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [19]),
        .Q(\I_0/hlctr_reg_n_0_[19] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[1] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [1]),
        .Q(\I_0/hlctr_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[20] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [20]),
        .Q(\I_0/hlctr_reg_n_0_[20] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[21] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [21]),
        .Q(\I_0/hlctr_reg_n_0_[21] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[22] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [22]),
        .Q(\I_0/hlctr_reg_n_0_[22] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[23] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [23]),
        .Q(\I_0/hlctr_reg_n_0_[23] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[24] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [24]),
        .Q(\I_0/hlctr_reg_n_0_[24] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[25] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [25]),
        .Q(\I_0/hlctr_reg_n_0_[25] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[26] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [26]),
        .Q(\I_0/hlctr_reg_n_0_[26] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[27] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [27]),
        .Q(\I_0/hlctr_reg_n_0_[27] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[28] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [28]),
        .Q(\I_0/hlctr_reg_n_0_[28] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[29] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [29]),
        .Q(\I_0/hlctr_reg_n_0_[29] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[2] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [2]),
        .Q(\I_0/hlctr_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[30] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [30]),
        .Q(\I_0/hlctr_reg_n_0_[30] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[31] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [31]),
        .Q(\I_0/hlctr_reg_n_0_[31] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[3] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [3]),
        .Q(\I_0/hlctr_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[4] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [4]),
        .Q(\I_0/hlctr_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[5] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [5]),
        .Q(\I_0/hlctr_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[6] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [6]),
        .Q(\I_0/hlctr_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[7] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [7]),
        .Q(\I_0/hlctr_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[8] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [8]),
        .Q(\I_0/hlctr_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/hlctr_reg[9] 
       (.C(clk15M),
        .CE(\I_0/hlctr0 ),
        .CLR(clear),
        .D(\I_0/hlctr [9]),
        .Q(\I_0/hlctr_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/i_austastung_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(i_austastung_i_1_n_0),
        .Q(\I_0/i_austastung ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_0/i_en_sync_last_reg 
       (.C(clk15M),
        .CE(reset),
        .D(\I_0/i_phase3 ),
        .Q(\I_0/i_en_sync_last ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_0/i_en_vertbr_last_reg 
       (.C(clk15M),
        .CE(reset),
        .D(\I_0/i_en_vertbr ),
        .Q(\I_0/i_en_vertbr_last ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/i_framereset_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(framereset_i_1_n_0),
        .Q(\I_0/i_framereset ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_phase4_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/i_phase4_inferred__0_carry_n_0 ,\I_0/i_phase4_inferred__0_carry_n_1 ,\I_0/i_phase4_inferred__0_carry_n_2 ,\I_0/i_phase4_inferred__0_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_phase4_inferred__0_carry_i_1_n_0,i_phase4_inferred__0_carry_i_2_n_0,i_phase4_inferred__0_carry_i_3_n_0,i_phase4_inferred__0_carry_i_4_n_0}),
        .S({i_phase4_inferred__0_carry_i_5_n_0,i_phase4_inferred__0_carry_i_6_n_0,i_phase4_inferred__0_carry_i_7_n_0,i_phase4_inferred__0_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_phase4_inferred__0_carry__0 
       (.CI(\I_0/i_phase4_inferred__0_carry_n_0 ),
        .CO({\I_0/i_phase4_inferred__0_carry__0_n_0 ,\I_0/i_phase4_inferred__0_carry__0_n_1 ,\I_0/i_phase4_inferred__0_carry__0_n_2 ,\I_0/i_phase4_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_phase4_inferred__0_carry__0_i_1_n_0,i_phase4_inferred__0_carry__0_i_2_n_0,i_phase4_inferred__0_carry__0_i_3_n_0,i_phase4_inferred__0_carry__0_i_4_n_0}),
        .S({i_phase4_inferred__0_carry__0_i_5_n_0,i_phase4_inferred__0_carry__0_i_6_n_0,i_phase4_inferred__0_carry__0_i_7_n_0,i_phase4_inferred__0_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_phase4_inferred__0_carry__1 
       (.CI(\I_0/i_phase4_inferred__0_carry__0_n_0 ),
        .CO({\I_0/i_phase4_inferred__0_carry__1_n_0 ,\I_0/i_phase4_inferred__0_carry__1_n_1 ,\I_0/i_phase4_inferred__0_carry__1_n_2 ,\I_0/i_phase4_inferred__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_phase4_inferred__0_carry__1_i_1_n_0,i_phase4_inferred__0_carry__1_i_2_n_0,i_phase4_inferred__0_carry__1_i_3_n_0,i_phase4_inferred__0_carry__1_i_4_n_0}),
        .S({i_phase4_inferred__0_carry__1_i_5_n_0,i_phase4_inferred__0_carry__1_i_6_n_0,i_phase4_inferred__0_carry__1_i_7_n_0,i_phase4_inferred__0_carry__1_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_phase4_inferred__0_carry__2 
       (.CI(\I_0/i_phase4_inferred__0_carry__1_n_0 ),
        .CO({\I_0/i_phase4 ,\I_0/i_phase4_inferred__0_carry__2_n_1 ,\I_0/i_phase4_inferred__0_carry__2_n_2 ,\I_0/i_phase4_inferred__0_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_phase4_inferred__0_carry__2_i_1_n_0,i_phase4_inferred__0_carry__2_i_2_n_0,i_phase4_inferred__0_carry__2_i_3_n_0,i_phase4_inferred__0_carry__2_i_4_n_0}),
        .S({i_phase4_inferred__0_carry__2_i_5_n_0,i_phase4_inferred__0_carry__2_i_6_n_0,i_phase4_inferred__0_carry__2_i_7_n_0,i_phase4_inferred__0_carry__2_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/i_phase_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(i_phase_i_1_n_0),
        .Q(phase));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/i_readmem_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(i_readmem_i_1_n_0),
        .Q(readmem));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_sync_c2_inferred__9_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/i_sync_c2_inferred__9_carry_n_0 ,\I_0/i_sync_c2_inferred__9_carry_n_1 ,\I_0/i_sync_c2_inferred__9_carry_n_2 ,\I_0/i_sync_c2_inferred__9_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_sync_c2_inferred__9_carry_i_1_n_0,i_sync_c2_inferred__9_carry_i_2_n_0,i_sync_c2_inferred__9_carry_i_3_n_0,i_sync_c2_inferred__9_carry_i_4_n_0}),
        .S({i_sync_c2_inferred__9_carry_i_5_n_0,i_sync_c2_inferred__9_carry_i_6_n_0,i_sync_c2_inferred__9_carry_i_7_n_0,i_sync_c2_inferred__9_carry_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_sync_c2_inferred__9_carry__0 
       (.CI(\I_0/i_sync_c2_inferred__9_carry_n_0 ),
        .CO({\I_0/i_sync_c2_inferred__9_carry__0_n_0 ,\I_0/i_sync_c2_inferred__9_carry__0_n_1 ,\I_0/i_sync_c2_inferred__9_carry__0_n_2 ,\I_0/i_sync_c2_inferred__9_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,i_sync_c2_inferred__9_carry__0_i_1_n_0}),
        .S({i_sync_c2_inferred__9_carry__0_i_2_n_0,i_sync_c2_inferred__9_carry__0_i_3_n_0,i_sync_c2_inferred__9_carry__0_i_4_n_0,i_sync_c2_inferred__9_carry__0_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_sync_c2_inferred__9_carry__1 
       (.CI(\I_0/i_sync_c2_inferred__9_carry__0_n_0 ),
        .CO({\I_0/i_sync_c2_inferred__9_carry__1_n_0 ,\I_0/i_sync_c2_inferred__9_carry__1_n_1 ,\I_0/i_sync_c2_inferred__9_carry__1_n_2 ,\I_0/i_sync_c2_inferred__9_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_sync_c2_inferred__9_carry__1_i_1_n_0,i_sync_c2_inferred__9_carry__1_i_2_n_0,i_sync_c2_inferred__9_carry__1_i_3_n_0,i_sync_c2_inferred__9_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/i_sync_c2_inferred__9_carry__2 
       (.CI(\I_0/i_sync_c2_inferred__9_carry__1_n_0 ),
        .CO({\I_0/i_sync_c223_in ,\I_0/i_sync_c2_inferred__9_carry__2_n_1 ,\I_0/i_sync_c2_inferred__9_carry__2_n_2 ,\I_0/i_sync_c2_inferred__9_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_sync_c2_inferred__9_carry__2_i_1_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_sync_c2_inferred__9_carry__2_i_2_n_0,i_sync_c2_inferred__9_carry__2_i_3_n_0,i_sync_c2_inferred__9_carry__2_i_4_n_0,i_sync_c2_inferred__9_carry__2_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_0/i_sync_c_reg[0] 
       (.C(clk15M),
        .CE(reset),
        .D(i_sync_c),
        .Q(\I_0/i_sync_c [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_0/i_sync_c_reg[1] 
       (.C(clk15M),
        .CE(reset),
        .D(\i_sync_c[1]_i_1_n_0 ),
        .Q(\I_0/i_sync_c [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr1_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/pixctr1_carry_n_0 ,\I_0/pixctr1_carry_n_1 ,\I_0/pixctr1_carry_n_2 ,\I_0/pixctr1_carry_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({pixctr1_carry_i_1_n_0,pixctr1_carry_i_2_n_0,pixctr1_carry_i_3_n_0,pixctr1_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr1_carry__0 
       (.CI(\I_0/pixctr1_carry_n_0 ),
        .CO({\I_0/pixctr1_carry__0_n_0 ,\I_0/pixctr1_carry__0_n_1 ,\I_0/pixctr1_carry__0_n_2 ,\I_0/pixctr1_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({pixctr1_carry__0_i_1_n_0,pixctr1_carry__0_i_2_n_0,pixctr1_carry__0_i_3_n_0,pixctr1_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr1_carry__1 
       (.CI(\I_0/pixctr1_carry__0_n_0 ),
        .CO({\I_0/pixctr1_carry__1_n_0 ,\I_0/pixctr1_carry__1_n_1 ,\I_0/pixctr1_carry__1_n_2 ,\I_0/pixctr1_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,pixctr1_carry__1_i_1_n_0,pixctr1_carry__1_i_2_n_0,pixctr1_carry__1_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_0/pixctr2_carry_n_0 ,\I_0/pixctr2_carry_n_1 ,\I_0/pixctr2_carry_n_2 ,\I_0/pixctr2_carry_n_3 }),
        .CYINIT(\I_0/pixctr_reg_n_0_ ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry_n_4 ,\I_0/pixctr2_carry_n_5 ,\I_0/pixctr2_carry_n_6 ,\I_0/pixctr2_carry_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[4] ,\I_0/pixctr_reg_n_0_[3] ,\I_0/pixctr_reg_n_0_[2] ,\I_0/pixctr_reg_n_0_[1] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__0 
       (.CI(\I_0/pixctr2_carry_n_0 ),
        .CO({\I_0/pixctr2_carry__0_n_0 ,\I_0/pixctr2_carry__0_n_1 ,\I_0/pixctr2_carry__0_n_2 ,\I_0/pixctr2_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__0_n_4 ,\I_0/pixctr2_carry__0_n_5 ,\I_0/pixctr2_carry__0_n_6 ,\I_0/pixctr2_carry__0_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[8] ,\I_0/pixctr_reg_n_0_[7] ,\I_0/pixctr_reg_n_0_[6] ,\I_0/pixctr_reg_n_0_[5] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__1 
       (.CI(\I_0/pixctr2_carry__0_n_0 ),
        .CO({\I_0/pixctr2_carry__1_n_0 ,\I_0/pixctr2_carry__1_n_1 ,\I_0/pixctr2_carry__1_n_2 ,\I_0/pixctr2_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__1_n_4 ,\I_0/pixctr2_carry__1_n_5 ,\I_0/pixctr2_carry__1_n_6 ,\I_0/pixctr2_carry__1_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[12] ,\I_0/pixctr_reg_n_0_[11] ,\I_0/pixctr_reg_n_0_[10] ,\I_0/pixctr_reg_n_0_[9] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__2 
       (.CI(\I_0/pixctr2_carry__1_n_0 ),
        .CO({\I_0/pixctr2_carry__2_n_0 ,\I_0/pixctr2_carry__2_n_1 ,\I_0/pixctr2_carry__2_n_2 ,\I_0/pixctr2_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__2_n_4 ,\I_0/pixctr2_carry__2_n_5 ,\I_0/pixctr2_carry__2_n_6 ,\I_0/pixctr2_carry__2_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[16] ,\I_0/pixctr_reg_n_0_[15] ,\I_0/pixctr_reg_n_0_[14] ,\I_0/pixctr_reg_n_0_[13] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__3 
       (.CI(\I_0/pixctr2_carry__2_n_0 ),
        .CO({\I_0/pixctr2_carry__3_n_0 ,\I_0/pixctr2_carry__3_n_1 ,\I_0/pixctr2_carry__3_n_2 ,\I_0/pixctr2_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__3_n_4 ,\I_0/pixctr2_carry__3_n_5 ,\I_0/pixctr2_carry__3_n_6 ,\I_0/pixctr2_carry__3_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[20] ,\I_0/pixctr_reg_n_0_[19] ,\I_0/pixctr_reg_n_0_[18] ,\I_0/pixctr_reg_n_0_[17] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__4 
       (.CI(\I_0/pixctr2_carry__3_n_0 ),
        .CO({\I_0/pixctr2_carry__4_n_0 ,\I_0/pixctr2_carry__4_n_1 ,\I_0/pixctr2_carry__4_n_2 ,\I_0/pixctr2_carry__4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__4_n_4 ,\I_0/pixctr2_carry__4_n_5 ,\I_0/pixctr2_carry__4_n_6 ,\I_0/pixctr2_carry__4_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[24] ,\I_0/pixctr_reg_n_0_[23] ,\I_0/pixctr_reg_n_0_[22] ,\I_0/pixctr_reg_n_0_[21] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__5 
       (.CI(\I_0/pixctr2_carry__4_n_0 ),
        .CO({\I_0/pixctr2_carry__5_n_0 ,\I_0/pixctr2_carry__5_n_1 ,\I_0/pixctr2_carry__5_n_2 ,\I_0/pixctr2_carry__5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__5_n_4 ,\I_0/pixctr2_carry__5_n_5 ,\I_0/pixctr2_carry__5_n_6 ,\I_0/pixctr2_carry__5_n_7 }),
        .S({\I_0/pixctr_reg_n_0_[28] ,\I_0/pixctr_reg_n_0_[27] ,\I_0/pixctr_reg_n_0_[26] ,\I_0/pixctr_reg_n_0_[25] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_0/pixctr2_carry__6 
       (.CI(\I_0/pixctr2_carry__5_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_0/pixctr2_carry__6_n_4 ,\I_0/pixctr2_carry__6_n_5 ,\I_0/pixctr2_carry__6_n_6 ,\I_0/pixctr2_carry__6_n_7 }),
        .S({\<const0>__0__0 ,\I_0/pixctr_reg_n_0_[31] ,\I_0/pixctr_reg_n_0_[30] ,\I_0/pixctr_reg_n_0_[29] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [0]),
        .Q(\I_0/pixctr_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [10]),
        .Q(\I_0/pixctr_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [11]),
        .Q(\I_0/pixctr_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[12] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [12]),
        .Q(\I_0/pixctr_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[13] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [13]),
        .Q(\I_0/pixctr_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[14] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [14]),
        .Q(\I_0/pixctr_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[15] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [15]),
        .Q(\I_0/pixctr_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[16] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [16]),
        .Q(\I_0/pixctr_reg_n_0_[16] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[17] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [17]),
        .Q(\I_0/pixctr_reg_n_0_[17] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[18] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [18]),
        .Q(\I_0/pixctr_reg_n_0_[18] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[19] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [19]),
        .Q(\I_0/pixctr_reg_n_0_[19] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [1]),
        .Q(\I_0/pixctr_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[20] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [20]),
        .Q(\I_0/pixctr_reg_n_0_[20] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[21] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [21]),
        .Q(\I_0/pixctr_reg_n_0_[21] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[22] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [22]),
        .Q(\I_0/pixctr_reg_n_0_[22] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[23] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [23]),
        .Q(\I_0/pixctr_reg_n_0_[23] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[24] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [24]),
        .Q(\I_0/pixctr_reg_n_0_[24] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[25] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [25]),
        .Q(\I_0/pixctr_reg_n_0_[25] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[26] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [26]),
        .Q(\I_0/pixctr_reg_n_0_[26] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[27] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [27]),
        .Q(\I_0/pixctr_reg_n_0_[27] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[28] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [28]),
        .Q(\I_0/pixctr_reg_n_0_[28] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[29] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [29]),
        .Q(\I_0/pixctr_reg_n_0_[29] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [2]),
        .Q(\I_0/pixctr_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[30] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [30]),
        .Q(\I_0/pixctr_reg_n_0_[30] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[31] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [31]),
        .Q(\I_0/pixctr_reg_n_0_[31] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [3]),
        .Q(\I_0/pixctr_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [4]),
        .Q(\I_0/pixctr_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [5]),
        .Q(\I_0/pixctr_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [6]),
        .Q(\I_0/pixctr_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [7]),
        .Q(\I_0/pixctr_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [8]),
        .Q(\I_0/pixctr_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/pixctr_reg[9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\I_0/pixctr [9]),
        .Q(\I_0/pixctr_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_0/sync_reg 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_0/p_1_in ),
        .Q(sync));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_1/abschnittu_reg[1] 
       (.C(clk),
        .CE(reset),
        .D(p_2_in),
        .Q(\I_1/abschnittu_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_10 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[4]),
        .O(\I_1/adr_reg_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_11 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[3]),
        .O(\I_1/adr_reg_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_12 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[2]),
        .O(\I_1/adr_reg_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_13 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[1]),
        .O(\I_1/adr_reg_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_14 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[0]),
        .O(\I_1/adr_reg_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_8 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[6]),
        .O(\I_1/adr_reg_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_1/adr_reg_i_9 
       (.I0(p_2_in__0[7]),
        .I1(p_2_in__0[5]),
        .O(\I_1/adr_reg_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[9]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[9]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[9]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[13]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[13]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[13]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[13]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[17]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[17]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[17]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[1]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[17]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[21]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[21]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[21]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[21]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[25]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[25]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[25]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[25]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[29]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[1]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[29]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[29]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[29]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[33]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[33]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[33]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[33]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[37]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[37]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[37]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[1]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[37]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[41]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[41]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[41]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[41]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[45]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[45]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[45]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[45]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[49]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[1]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[49]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[49]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[49]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[53]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[53]_i_1_n_6 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[53]_i_1_n_5 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[53]_i_1_n_4 ),
        .PRE(i_phase_i_2_n_0),
        .Q(\I_1/ctr90_48_reg [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[57]_i_1_n_7 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[57]_i_1_n_6 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[57]_i_1_n_5 ),
        .PRE(i_phase_i_2_n_0),
        .Q(\I_1/ctr90_48_reg [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[5]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[57]_i_1_n_4 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr90_48_reg[61]_i_1_n_7 ),
        .PRE(pixctr),
        .Q(\I_1/ctr90_48_reg [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[61]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr90_48_reg[61]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[5]_i_1_n_6 ),
        .Q(\I_1/ctr90_48_reg [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[5]_i_1_n_5 ),
        .Q(\I_1/ctr90_48_reg [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[5]_i_1_n_4 ),
        .Q(\I_1/ctr90_48_reg [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr90_48_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\ctr90_48_reg[9]_i_1_n_7 ),
        .Q(\I_1/ctr90_48_reg [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[9]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[9]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[9]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[13]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[13]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[13]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[13]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[17]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[17]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[17]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[1]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[17]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[21]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[21]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[21]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[21]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[25]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[25]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[25]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[25]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[29]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[1]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[29]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[29]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[32] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[29]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[33] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[33]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[34] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[33]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[35] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[33]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[36] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[33]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[37] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[37]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[38] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[37]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[39] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[37]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[1]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[40] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[37]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[41] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[41]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[42] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[41]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[43] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[41]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[44] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[41]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[45] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[45]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[46] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[45]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[47] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[45]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[48] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[45]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[49] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[49]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[1]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[50] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[49]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[51] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[49]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[52] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[49]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[53] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[53]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[54] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[53]_i_1_n_6 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[55] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[53]_i_1_n_5 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[56] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[53]_i_1_n_4 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[57] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[57]_i_1_n_7 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[58] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[57]_i_1_n_6 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[59] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[57]_i_1_n_5 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[5]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[60] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[57]_i_1_n_4 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[61] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[61]_i_1_n_7 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[62] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[61]_i_1_n_6 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDPE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_PRE_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\ctr_48_reg[61]_i_1_n_5 ),
        .PRE(pixctr),
        .Q(\I_1/ctr_48_reg [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[5]_i_1_n_6 ),
        .Q(\I_1/ctr_48_reg [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[5]_i_1_n_5 ),
        .Q(\I_1/ctr_48_reg [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[5]_i_1_n_4 ),
        .Q(\I_1/ctr_48_reg [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/ctr_48_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(pixctr),
        .D(\ctr_48_reg[9]_i_1_n_7 ),
        .Q(\I_1/ctr_48_reg [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[10]_i_1 
       (.I0(\data_reg[12]_i_2__0_n_6 ),
        .I1(\I_2/adr_reg_n_21 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[11]_i_1 
       (.I0(\data_reg[12]_i_2__0_n_5 ),
        .I1(\I_2/adr_reg_n_20 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[12]_i_1 
       (.I0(\data_reg[12]_i_2__0_n_4 ),
        .I1(\I_2/adr_reg_n_19 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[12]_i_3 
       (.I0(\I_2/adr_reg_n_19 ),
        .O(\I_1/data[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[12]_i_4 
       (.I0(\I_2/adr_reg_n_20 ),
        .O(\I_1/data[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[12]_i_5 
       (.I0(\I_2/adr_reg_n_21 ),
        .O(\I_1/data[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[12]_i_6 
       (.I0(\I_2/adr_reg_n_22 ),
        .O(\I_1/data[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[13]_i_1 
       (.I0(\data_reg[15]_i_2__0_n_7 ),
        .I1(\I_2/adr_reg_n_18 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[14]_i_1 
       (.I0(\data_reg[15]_i_2__0_n_6 ),
        .I1(\I_2/adr_reg_n_17 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \I_1/data[15]_i_1 
       (.I0(\I_1/abschnittu_reg_n_0_ ),
        .I1(\data_reg[15]_i_2__0_n_1 ),
        .O(\I_1/data[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[15]_i_3 
       (.I0(\I_2/adr_reg_n_17 ),
        .O(\I_1/data[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[15]_i_4 
       (.I0(\I_2/adr_reg_n_18 ),
        .O(\I_1/data[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[1]_i_1 
       (.I0(\data_reg[4]_i_2__0_n_7 ),
        .I1(\I_2/adr_reg_n_30 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[2]_i_1 
       (.I0(\data_reg[4]_i_2__0_n_6 ),
        .I1(\I_2/adr_reg_n_29 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[3]_i_1 
       (.I0(\data_reg[4]_i_2__0_n_5 ),
        .I1(\I_2/adr_reg_n_28 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[4]_i_1 
       (.I0(\data_reg[4]_i_2__0_n_4 ),
        .I1(\I_2/adr_reg_n_27 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[4]_i_3 
       (.I0(\I_2/adr_reg_n_31 ),
        .O(\I_1/data[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[4]_i_4 
       (.I0(\I_2/adr_reg_n_27 ),
        .O(\I_1/data[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[4]_i_5 
       (.I0(\I_2/adr_reg_n_28 ),
        .O(\I_1/data[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[4]_i_6 
       (.I0(\I_2/adr_reg_n_29 ),
        .O(\I_1/data[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[4]_i_7 
       (.I0(\I_2/adr_reg_n_30 ),
        .O(\I_1/data[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[5]_i_1 
       (.I0(\data_reg[8]_i_2__0_n_7 ),
        .I1(\I_2/adr_reg_n_26 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[6]_i_1 
       (.I0(\data_reg[8]_i_2__0_n_6 ),
        .I1(\I_2/adr_reg_n_25 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[7]_i_1 
       (.I0(\data_reg[8]_i_2__0_n_5 ),
        .I1(\I_2/adr_reg_n_24 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[8]_i_1 
       (.I0(\data_reg[8]_i_2__0_n_4 ),
        .I1(\I_2/adr_reg_n_23 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[8]_i_3 
       (.I0(\I_2/adr_reg_n_23 ),
        .O(\I_1/data[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[8]_i_4 
       (.I0(\I_2/adr_reg_n_24 ),
        .O(\I_1/data[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[8]_i_5 
       (.I0(\I_2/adr_reg_n_25 ),
        .O(\I_1/data[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_1/data[8]_i_6 
       (.I0(\I_2/adr_reg_n_26 ),
        .O(\I_1/data[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_1/data[9]_i_1 
       (.I0(\data_reg[12]_i_2__0_n_7 ),
        .I1(\I_2/adr_reg_n_22 ),
        .I2(\I_1/abschnittu_reg_n_0_ ),
        .O(\I_1/data[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_2/adr_reg_n_31 ),
        .Q(\I_1/data_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data ),
        .Q(\I_1/data_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[11]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[12]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[12] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[13]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[13] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[14]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[14] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[15]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[15] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[1]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[2]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[3]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[4]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[5]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[6]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[7]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[8]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_1/data_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_1/data[9]_i_1_n_0 ),
        .Q(\I_1/data_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_2/abschnittu_reg[1] 
       (.C(clk),
        .CE(reset),
        .D(p_3_in),
        .Q(abschnittu),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}}" *) 
  (* RTL_RAM_BITS = "1920" *) 
  (* RTL_RAM_NAME = "I_2/adr" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h183316A7151B138E120010720EE30D530BC30A3208A10710057E03ED025B00C9),
    .INIT_01(256'h30412ECC2D542BDB2A6128E5276725E7246722E421611FDC1E561CCF1B4619BD),
    .INIT_02(256'h4674452343D0427941203FC53E673D073BA43A3F38D8376F36033496332631B4),
    .INIT_03(256'h59F358D357B05689555F5432530151CE50974F5D4E204CE04B9D4A57490E47C3),
    .INIT_04(256'h69FC69196831674566566562646B63706271616E60675F5D5E4F5D3D5C285B0F),
    .INIT_05(256'h75F3755474B1740A735E72AE71F9714070826FC06EFA6E306D616C8E6BB76ADB),
    .INIT_06(256'h7D617D0E7CB67C597BF77B917B257AB57A4179C7794978C6783F77B37722768D),
    .INIT_07(256'h7FFE7FF97FEF7FE07FCD7FB47F967F747F4C7F207EEF7EB97E7E7E3E7DF97DB0),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("PERFORMANCE"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("WRITE_FIRST"),
    .WRITE_MODE_B("WRITE_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(0)) 
    \I_2/adr_reg 
       (.ADDRARDADDR({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_2/adr_reg_i_1_n_0 ,\I_2/adr_reg_i_2_n_0 ,\I_2/adr_reg_i_3_n_0 ,\I_2/adr_reg_i_4_n_0 ,\I_2/adr_reg_i_5_n_0 ,\I_2/adr_reg_i_6_n_0 ,\I_2/adr_reg_i_7_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ADDRBWRADDR({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/adr_reg_i_8_n_0 ,\I_1/adr_reg_i_9_n_0 ,\I_1/adr_reg_i_10_n_0 ,\I_1/adr_reg_i_11_n_0 ,\I_1/adr_reg_i_12_n_0 ,\I_1/adr_reg_i_13_n_0 ,\I_1/adr_reg_i_14_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIBDI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const1>__0__0 ,\<const1>__0__0 }),
        .DOADO({\I_2/adr_reg_n_0 ,\I_2/adr_reg_n_1 ,\I_2/adr_reg_n_2 ,\I_2/adr_reg_n_3 ,\I_2/adr_reg_n_4 ,\I_2/adr_reg_n_5 ,\I_2/adr_reg_n_6 ,\I_2/adr_reg_n_7 ,\I_2/adr_reg_n_8 ,\I_2/adr_reg_n_9 ,\I_2/adr_reg_n_10 ,\I_2/adr_reg_n_11 ,\I_2/adr_reg_n_12 ,\I_2/adr_reg_n_13 ,\I_2/adr_reg_n_14 ,p_1_in[0]}),
        .DOBDO({\I_2/adr_reg_n_16 ,\I_2/adr_reg_n_17 ,\I_2/adr_reg_n_18 ,\I_2/adr_reg_n_19 ,\I_2/adr_reg_n_20 ,\I_2/adr_reg_n_21 ,\I_2/adr_reg_n_22 ,\I_2/adr_reg_n_23 ,\I_2/adr_reg_n_24 ,\I_2/adr_reg_n_25 ,\I_2/adr_reg_n_26 ,\I_2/adr_reg_n_27 ,\I_2/adr_reg_n_28 ,\I_2/adr_reg_n_29 ,\I_2/adr_reg_n_30 ,\I_2/adr_reg_n_31 }),
        .ENARDEN(reset),
        .ENBWREN(reset),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\<const0>__0__0 ,\<const0>__0__0 }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_1 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[6]),
        .O(\I_2/adr_reg_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_2 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[5]),
        .O(\I_2/adr_reg_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_3 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[4]),
        .O(\I_2/adr_reg_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_4 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[3]),
        .O(\I_2/adr_reg_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_5 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[2]),
        .O(\I_2/adr_reg_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_6 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[1]),
        .O(\I_2/adr_reg_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_2/adr_reg_i_7 
       (.I0(p_3_in__0[7]),
        .I1(p_3_in__0[0]),
        .O(\I_2/adr_reg_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[10]_i_1 
       (.I0(data0[10]),
        .I1(\I_2/adr_reg_n_5 ),
        .I2(abschnittu),
        .O(p_1_in[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[11]_i_1 
       (.I0(data0[11]),
        .I1(\I_2/adr_reg_n_4 ),
        .I2(abschnittu),
        .O(p_1_in[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[12]_i_1 
       (.I0(data0[12]),
        .I1(\I_2/adr_reg_n_3 ),
        .I2(abschnittu),
        .O(p_1_in[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[12]_i_3 
       (.I0(\I_2/adr_reg_n_3 ),
        .O(\I_2/data ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[12]_i_4 
       (.I0(\I_2/adr_reg_n_4 ),
        .O(\I_2/data[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[12]_i_5 
       (.I0(\I_2/adr_reg_n_5 ),
        .O(\I_2/data[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[12]_i_6 
       (.I0(\I_2/adr_reg_n_6 ),
        .O(\I_2/data[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[13]_i_1 
       (.I0(data0[13]),
        .I1(\I_2/adr_reg_n_2 ),
        .I2(abschnittu),
        .O(p_1_in[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[14]_i_1 
       (.I0(data0[14]),
        .I1(\I_2/adr_reg_n_1 ),
        .I2(abschnittu),
        .O(p_1_in[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \I_2/data[15]_i_1 
       (.I0(abschnittu),
        .I1(\data_reg[15]_i_2_n_1 ),
        .O(p_1_in[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[15]_i_3 
       (.I0(\I_2/adr_reg_n_1 ),
        .O(\I_2/data[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[15]_i_4 
       (.I0(\I_2/adr_reg_n_2 ),
        .O(\I_2/data[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[1]_i_1 
       (.I0(data0[1]),
        .I1(\I_2/adr_reg_n_14 ),
        .I2(abschnittu),
        .O(p_1_in[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[2]_i_1 
       (.I0(data0[2]),
        .I1(\I_2/adr_reg_n_13 ),
        .I2(abschnittu),
        .O(p_1_in[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[3]_i_1 
       (.I0(data0[3]),
        .I1(\I_2/adr_reg_n_12 ),
        .I2(abschnittu),
        .O(p_1_in[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[4]_i_1 
       (.I0(data0[4]),
        .I1(\I_2/adr_reg_n_11 ),
        .I2(abschnittu),
        .O(p_1_in[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[4]_i_3 
       (.I0(p_1_in[0]),
        .O(\I_2/data[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[4]_i_4 
       (.I0(\I_2/adr_reg_n_11 ),
        .O(\I_2/data[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[4]_i_5 
       (.I0(\I_2/adr_reg_n_12 ),
        .O(\I_2/data[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[4]_i_6 
       (.I0(\I_2/adr_reg_n_13 ),
        .O(\I_2/data[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[4]_i_7 
       (.I0(\I_2/adr_reg_n_14 ),
        .O(\I_2/data[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[5]_i_1 
       (.I0(data0[5]),
        .I1(\I_2/adr_reg_n_10 ),
        .I2(abschnittu),
        .O(p_1_in[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[6]_i_1 
       (.I0(data0[6]),
        .I1(\I_2/adr_reg_n_9 ),
        .I2(abschnittu),
        .O(p_1_in[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[7]_i_1 
       (.I0(data0[7]),
        .I1(\I_2/adr_reg_n_8 ),
        .I2(abschnittu),
        .O(p_1_in[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[8]_i_1 
       (.I0(data0[8]),
        .I1(\I_2/adr_reg_n_7 ),
        .I2(abschnittu),
        .O(p_1_in[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[8]_i_3 
       (.I0(\I_2/adr_reg_n_7 ),
        .O(\I_2/data[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[8]_i_4 
       (.I0(\I_2/adr_reg_n_8 ),
        .O(\I_2/data[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[8]_i_5 
       (.I0(\I_2/adr_reg_n_9 ),
        .O(\I_2/data[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_2/data[8]_i_6 
       (.I0(\I_2/adr_reg_n_10 ),
        .O(\I_2/data[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \I_2/data[9]_i_1 
       (.I0(data0[9]),
        .I1(\I_2/adr_reg_n_6 ),
        .I2(abschnittu),
        .O(p_1_in[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[0]),
        .Q(data[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[10]),
        .Q(data[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[11]),
        .Q(data[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[12]),
        .Q(data[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[13]),
        .Q(data[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[14]),
        .Q(data[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[15]),
        .Q(data[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[1]),
        .Q(data[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[2]),
        .Q(data[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[3]),
        .Q(data[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[4]),
        .Q(data[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[5]),
        .Q(data[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[6]),
        .Q(data[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[7]),
        .Q(data[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[8]),
        .Q(data[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_2/data_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(p_1_in[9]),
        .Q(data[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_3/minusOp_carry_n_0 ,\I_3/minusOp_carry_n_1 ,\I_3/minusOp_carry_n_2 ,\I_3/minusOp_carry_n_3 }),
        .CYINIT(\I_3/minusOp_inferred__0__0_i_2_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_3/minusOp_carry_n_4 ,\I_3/minusOp_carry_n_5 ,\I_3/minusOp_carry_n_6 ,\I_3/minusOp_carry_n_7 }),
        .S({\I_3/minusOp_carry_i_1_n_0 ,\I_3/minusOp_carry_i_2_n_0 ,\I_3/minusOp_carry_i_3_n_0 ,\I_3/minusOp_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_carry__0 
       (.CI(\I_3/minusOp_carry_n_0 ),
        .CO({\I_3/minusOp_carry__0_n_0 ,\I_3/minusOp_carry__0_n_1 ,\I_3/minusOp_carry__0_n_2 ,\I_3/minusOp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(in_r[3:0]),
        .O({\I_3/minusOp_carry__0_n_4 ,\I_3/minusOp_carry__0_n_5 ,\I_3/minusOp_carry__0_n_6 ,\I_3/minusOp_carry__0_n_7 }),
        .S({minusOp_carry__0_i_1_n_0,minusOp_carry__0_i_2_n_0,minusOp_carry__0_i_3_n_0,minusOp_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_carry__1 
       (.CI(\I_3/minusOp_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,in_r[4]}),
        .O({\I_3/minusOp_carry__1_n_4 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_6 ,\I_3/minusOp_carry__1_n_7 }),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\I_3/plusOp__0_carry__1_n_5 ,minusOp_carry__1_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_carry_i_1 
       (.I0(plusOp18[4]),
        .O(\I_3/minusOp_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_carry_i_2 
       (.I0(plusOp18[3]),
        .O(\I_3/minusOp_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_carry_i_3 
       (.I0(plusOp18[2]),
        .O(\I_3/minusOp_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_carry_i_4 
       (.I0(plusOp18[1]),
        .O(\I_3/minusOp_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* XILINX_LEGACY_PRIM = "(MUXCY,XORCY)" *) 
  CARRY4 \I_3/minusOp_inferred__0__0_CARRY4 
       (.CI(lopt),
        .CYINIT(\I_3/minusOp_inferred__0__0_i_2_n_0 ),
        .O({\I_3/minusOp_inferred__0__0_CARRY4_n_4 ,\I_3/minusOp_inferred__0__0_CARRY4_n_5 ,\I_3/minusOp_inferred__0__0_CARRY4_n_6 ,\I_3/minusOp_inferred__0__0_n_0 }),
        .S(\I_3/minusOp_inferred__0__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND \I_3/minusOp_inferred__0__0_CARRY4_GND 
       (.G(lopt));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0__0_i_1 
       (.I0(plusOp18[1]),
        .O(\I_3/minusOp_inferred__0__0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0__0_i_2 
       (.I0(plusOp18[0]),
        .O(\I_3/minusOp_inferred__0__0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_inferred__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_3/minusOp_inferred__0_carry_n_0 ,\I_3/minusOp_inferred__0_carry_n_1 ,\I_3/minusOp_inferred__0_carry_n_2 ,\I_3/minusOp_inferred__0_carry_n_3 }),
        .CYINIT(\I_3/minusOp_inferred__0__0_i_2_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_3/minusOp_inferred__0_carry_n_4 ,\I_3/minusOp_inferred__0_carry_n_5 ,\I_3/minusOp_inferred__0_carry_n_6 ,\I_3/minusOp_inferred__0_carry_n_7 }),
        .S({\I_3/minusOp_inferred__0_carry_i_1_n_0 ,\I_3/minusOp_inferred__0_carry_i_2_n_0 ,\I_3/minusOp_inferred__0_carry_i_3_n_0 ,\I_3/minusOp_inferred__0_carry_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_inferred__0_carry__0 
       (.CI(\I_3/minusOp_inferred__0_carry_n_0 ),
        .CO({\I_3/minusOp_inferred__0_carry__0_n_0 ,\I_3/minusOp_inferred__0_carry__0_n_1 ,\I_3/minusOp_inferred__0_carry__0_n_2 ,\I_3/minusOp_inferred__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(in_b[3:0]),
        .O({\I_3/minusOp_inferred__0_carry__0_n_4 ,\I_3/minusOp_inferred__0_carry__0_n_5 ,\I_3/minusOp_inferred__0_carry__0_n_6 ,\I_3/minusOp_inferred__0_carry__0_n_7 }),
        .S({minusOp_inferred__0_carry__0_i_1_n_0,minusOp_inferred__0_carry__0_i_2_n_0,minusOp_inferred__0_carry__0_i_3_n_0,minusOp_inferred__0_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/minusOp_inferred__0_carry__1 
       (.CI(\I_3/minusOp_inferred__0_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,in_b[4]}),
        .O({\I_3/minusOp_inferred__0_carry__1_n_4 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_6 ,\I_3/minusOp_inferred__0_carry__1_n_7 }),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\I_3/plusOp__0_carry__1_n_5 ,minusOp_inferred__0_carry__1_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0_carry_i_1 
       (.I0(plusOp18[4]),
        .O(\I_3/minusOp_inferred__0_carry_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0_carry_i_2 
       (.I0(plusOp18[3]),
        .O(\I_3/minusOp_inferred__0_carry_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0_carry_i_3 
       (.I0(plusOp18[2]),
        .O(\I_3/minusOp_inferred__0_carry_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \I_3/minusOp_inferred__0_carry_i_4 
       (.I0(plusOp18[1]),
        .O(\I_3/minusOp_inferred__0_carry_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_3/multOp 
       (.A({\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_5 ,\I_3/minusOp_carry__1_n_6 ,\I_3/minusOp_carry__1_n_7 ,\I_3/minusOp_carry__0_n_4 ,\I_3/minusOp_carry__0_n_5 ,\I_3/minusOp_carry__0_n_6 ,\I_3/minusOp_carry__0_n_7 ,\I_3/minusOp_carry_n_4 ,\I_3/minusOp_carry_n_5 ,\I_3/minusOp_carry_n_6 ,\I_3/minusOp_carry_n_7 ,plusOp18[0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk15M),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\I_3/multOp_n_58 ,\I_3/multOp_n_59 ,\I_3/multOp_n_60 ,\I_3/multOp_n_61 ,\I_3/multOp_n_62 ,\I_3/multOp_n_63 ,\I_3/multOp_n_64 ,\I_3/multOp_n_65 ,\I_3/multOp_n_66 ,\I_3/multOp_n_67 ,\I_3/multOp_n_68 ,\I_3/multOp_n_69 ,\I_3/multOp_n_70 ,\I_3/multOp_n_71 ,\I_3/multOp_n_72 ,\I_3/multOp_n_73 ,\I_3/multOp_n_74 ,\I_3/multOp_n_75 ,\I_3/multOp_n_76 ,\I_3/multOp_n_77 ,\I_3/multOp_n_78 ,\I_3/multOp_n_79 ,\I_3/multOp_n_80 ,\I_3/multOp_n_81 ,\I_3/multOp_n_82 ,\I_3/multOp_n_83 ,\I_3/multOp_n_84 ,\I_3/multOp_n_85 ,\I_3/multOp_n_86 ,\I_3/multOp_n_87 ,\I_3/multOp_n_88 ,\I_3/multOp_n_89 ,\I_3/multOp_n_90 ,\I_3/multOp_n_91 ,\I_3/multOp_n_92 ,\I_3/multOp_n_93 ,\I_3/multOp_n_94 ,\I_3/multOp_n_95 ,\I_3/multOp_n_96 ,\I_3/multOp_n_97 ,\I_3/multOp_n_98 ,\I_3/multOp_n_99 ,\I_3/multOp_n_100 ,\I_3/multOp_n_101 ,\I_3/multOp_n_102 ,\I_3/multOp_n_103 ,\I_3/multOp_n_104 ,\I_3/multOp_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(1),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_3/multOp__0 
       (.A({\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_5 ,\I_3/minusOp_inferred__0_carry__1_n_6 ,\I_3/minusOp_inferred__0_carry__1_n_7 ,\I_3/minusOp_inferred__0_carry__0_n_4 ,\I_3/minusOp_inferred__0_carry__0_n_5 ,\I_3/minusOp_inferred__0_carry__0_n_6 ,\I_3/minusOp_inferred__0_carry__0_n_7 ,\I_3/minusOp_inferred__0_carry_n_4 ,\I_3/minusOp_inferred__0_carry_n_5 ,\I_3/minusOp_inferred__0_carry_n_6 ,\I_3/minusOp_inferred__0__0_n_0 ,plusOp18[0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const1>__0__0 ),
        .CLK(clk15M),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\I_3/multOp__0_n_58 ,\I_3/multOp__0_n_59 ,\I_3/multOp__0_n_60 ,\I_3/multOp__0_n_61 ,\I_3/multOp__0_n_62 ,\I_3/multOp__0_n_63 ,\I_3/multOp__0_n_64 ,\I_3/multOp__0_n_65 ,\I_3/multOp__0_n_66 ,\I_3/multOp__0_n_67 ,\I_3/multOp__0_n_68 ,\I_3/multOp__0_n_69 ,\I_3/multOp__0_n_70 ,\I_3/multOp__0_n_71 ,\I_3/multOp__0_n_72 ,\I_3/multOp__0_n_73 ,\I_3/multOp__0_n_74 ,\I_3/multOp__0_n_75 ,\I_3/multOp__0_n_76 ,\I_3/multOp__0_n_77 ,\I_3/multOp__0_n_78 ,\I_3/multOp__0_n_79 ,\I_3/multOp__0_n_80 ,\I_3/multOp__0_n_81 ,\I_3/multOp__0_n_82 ,\I_3/multOp__0_n_83 ,\I_3/multOp__0_n_84 ,\I_3/multOp__0_n_85 ,\I_3/multOp__0_n_86 ,\I_3/multOp__0_n_87 ,\I_3/multOp__0_n_88 ,\I_3/multOp__0_n_89 ,\I_3/multOp__0_n_90 ,\I_3/multOp__0_n_91 ,\I_3/multOp__0_n_92 ,\I_3/multOp__0_n_93 ,\I_3/multOp__0_n_94 ,\I_3/multOp__0_n_95 ,\I_3/multOp__0_n_96 ,\I_3/multOp__0_n_97 ,\I_3/multOp__0_n_98 ,\I_3/multOp__0_n_99 ,\I_3/multOp__0_n_100 ,\I_3/multOp__0_n_101 ,\I_3/multOp__0_n_102 ,\I_3/multOp__0_n_103 ,\I_3/multOp__0_n_104 ,\I_3/multOp__0_n_105 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_3/out_y_reg_c 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\<const1>__0__0 ),
        .Q(\I_3/out_y_reg_c_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/plusOp__0_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_3/plusOp__0_carry_n_0 ,\I_3/plusOp__0_carry_n_1 ,\I_3/plusOp__0_carry_n_2 ,\I_3/plusOp__0_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({plusOp__0_carry_i_1_n_0,plusOp__0_carry_i_2_n_0,g0_b0__0_n_0,\<const0>__0__0 }),
        .O(plusOp18[3:0]),
        .S({plusOp__0_carry_i_3_n_0,plusOp__0_carry_i_4_n_0,plusOp__0_carry_i_5_n_0,g0_b0__0__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/plusOp__0_carry__0 
       (.CI(\I_3/plusOp__0_carry_n_0 ),
        .CO({\I_3/plusOp__0_carry__0_n_0 ,\I_3/plusOp__0_carry__0_n_1 ,\I_3/plusOp__0_carry__0_n_2 ,\I_3/plusOp__0_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({plusOp__0_carry__0_i_1_n_0,plusOp__0_carry__0_i_2_n_0,plusOp__0_carry__0_i_3_n_0,plusOp__0_carry__0_i_4_n_0}),
        .O(plusOp18[7:4]),
        .S({plusOp__0_carry__0_i_5_n_0,plusOp__0_carry__0_i_6_n_0,plusOp__0_carry__0_i_7_n_0,plusOp__0_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_3/plusOp__0_carry__1 
       (.CI(\I_3/plusOp__0_carry__0_n_0 ),
        .CO({\I_3/plusOp__0_carry__1_n_0 ,\I_3/plusOp__0_carry__1_n_1 ,plusOp18[10],\I_3/plusOp__0_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,g0_b9_n_0,plusOp__0_carry__1_i_1_n_0}),
        .O({\I_3/plusOp__0_carry__1_n_4 ,\I_3/plusOp__0_carry__1_n_5 ,plusOp18[9:8]}),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,g0_b9__0_n_0,plusOp__0_carry__1_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/multOp 
       (.A({\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_5 ,\I_4/multOp_i_1_n_6 ,\I_4/multOp_i_1_n_7 ,\I_4/multOp_i_2_n_4 ,\I_4/multOp_i_2_n_5 ,\I_4/multOp_i_2_n_6 ,\I_4/multOp_i_2_n_7 ,\I_4/multOp_i_3_n_4 ,\I_4/multOp_i_3_n_5 ,\I_4/multOp_i_3_n_6 ,\I_4/multOp_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\I_4/multOp_n_106 ,\I_4/multOp_n_107 ,\I_4/multOp_n_108 ,\I_4/multOp_n_109 ,\I_4/multOp_n_110 ,\I_4/multOp_n_111 ,\I_4/multOp_n_112 ,\I_4/multOp_n_113 ,\I_4/multOp_n_114 ,\I_4/multOp_n_115 ,\I_4/multOp_n_116 ,\I_4/multOp_n_117 ,\I_4/multOp_n_118 ,\I_4/multOp_n_119 ,\I_4/multOp_n_120 ,\I_4/multOp_n_121 ,\I_4/multOp_n_122 ,\I_4/multOp_n_123 ,\I_4/multOp_n_124 ,\I_4/multOp_n_125 ,\I_4/multOp_n_126 ,\I_4/multOp_n_127 ,\I_4/multOp_n_128 ,\I_4/multOp_n_129 ,\I_4/multOp_n_130 ,\I_4/multOp_n_131 ,\I_4/multOp_n_132 ,\I_4/multOp_n_133 ,\I_4/multOp_n_134 ,\I_4/multOp_n_135 ,\I_4/multOp_n_136 ,\I_4/multOp_n_137 ,\I_4/multOp_n_138 ,\I_4/multOp_n_139 ,\I_4/multOp_n_140 ,\I_4/multOp_n_141 ,\I_4/multOp_n_142 ,\I_4/multOp_n_143 ,\I_4/multOp_n_144 ,\I_4/multOp_n_145 ,\I_4/multOp_n_146 ,\I_4/multOp_n_147 ,\I_4/multOp_n_148 ,\I_4/multOp_n_149 ,\I_4/multOp_n_150 ,\I_4/multOp_n_151 ,\I_4/multOp_n_152 ,\I_4/multOp_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp__39_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/multOp__39_carry_n_0 ,\I_4/multOp__39_carry_n_1 ,\I_4/multOp__39_carry_n_2 ,\I_4/multOp__39_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry_i_1__0_n_0,multOp__39_carry_i_2__0_n_0,multOp__39_carry_i_3__0_n_0,\<const0>__0__0 }),
        .O(multOp0[6:3]),
        .S({multOp__39_carry_i_4__0_n_0,multOp__39_carry_i_5__0_n_0,multOp__39_carry_i_6__0_n_0,multOp__39_carry_i_7__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp__39_carry__0 
       (.CI(\I_4/multOp__39_carry_n_0 ),
        .CO({\I_4/multOp__39_carry__0_n_0 ,\I_4/multOp__39_carry__0_n_1 ,\I_4/multOp__39_carry__0_n_2 ,\I_4/multOp__39_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry__0_i_1__0_n_0,multOp__39_carry__0_i_2__0_n_0,multOp__39_carry__0_i_3__0_n_0,multOp__39_carry__0_i_4__0_n_0}),
        .O(multOp0[10:7]),
        .S({multOp__39_carry__0_i_5__0_n_0,multOp__39_carry__0_i_6__0_n_0,multOp__39_carry__0_i_7__0_n_0,multOp__39_carry__0_i_8__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp__39_carry__1 
       (.CI(\I_4/multOp__39_carry__0_n_0 ),
        .CO({\I_4/multOp__39_carry__1_n_0 ,\I_4/multOp__39_carry__1_n_1 ,\I_4/multOp__39_carry__1_n_2 ,\I_4/multOp__39_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry__1_i_1__0_n_0,multOp__39_carry__1_i_2__0_n_0,multOp__39_carry__1_i_3__0_n_0,multOp__39_carry__1_i_4__0_n_0}),
        .O(multOp0[14:11]),
        .S({multOp__39_carry__1_i_5__0_n_0,multOp__39_carry__1_i_6__0_n_0,multOp__39_carry__1_i_7__0_n_0,multOp__39_carry__1_i_8__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp__39_carry__2 
       (.CI(\I_4/multOp__39_carry__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_4/multOp__39_carry__2_n_4 ,\I_4/multOp__39_carry__2_n_5 ,\I_4/multOp__39_carry__2_n_6 ,multOp0[15]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,multOp__39_carry__2_i_1__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/multOp_carry_n_0 ,\I_4/multOp_carry_n_1 ,\I_4/multOp_carry_n_2 ,\I_4/multOp_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/plusOp_inferred__6_carry_n_6 ,\I_4/plusOp_inferred__6_carry_n_7 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\I_4/multOp_carry_n_4 ,multOp0[2:0]}),
        .S({multOp_carry_i_1__0_n_0,multOp_carry_i_2__0_n_0,multOp_carry_i_3__0_n_0,\I_4/plusOp_inferred__6_carry_n_7 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_carry__0 
       (.CI(\I_4/multOp_carry_n_0 ),
        .CO({\I_4/multOp_carry__0_n_0 ,\I_4/multOp_carry__0_n_1 ,\I_4/multOp_carry__0_n_2 ,\I_4/multOp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/plusOp_inferred__6_carry__0_n_6 ,\I_4/plusOp_inferred__6_carry__0_n_7 ,\I_4/plusOp_inferred__6_carry_n_4 ,\I_4/plusOp_inferred__6_carry_n_5 }),
        .O({\I_4/multOp_carry__0_n_4 ,\I_4/multOp_carry__0_n_5 ,\I_4/multOp_carry__0_n_6 ,\I_4/multOp_carry__0_n_7 }),
        .S({multOp_carry__0_i_1__0_n_0,multOp_carry__0_i_2__0_n_0,multOp_carry__0_i_3__0_n_0,multOp_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_carry__1 
       (.CI(\I_4/multOp_carry__0_n_0 ),
        .CO({\I_4/multOp_carry__1_n_0 ,\I_4/multOp_carry__1_n_1 ,\I_4/multOp_carry__1_n_2 ,\I_4/multOp_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/plusOp_inferred__6_carry__1_n_6 ,\I_4/plusOp_inferred__6_carry__1_n_7 ,\I_4/plusOp_inferred__6_carry__0_n_4 ,\I_4/plusOp_inferred__6_carry__0_n_5 }),
        .O({\I_4/multOp_carry__1_n_4 ,\I_4/multOp_carry__1_n_5 ,\I_4/multOp_carry__1_n_6 ,\I_4/multOp_carry__1_n_7 }),
        .S({multOp_carry__1_i_1__0_n_0,multOp_carry__1_i_2__0_n_0,multOp_carry__1_i_3__0_n_0,multOp_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_carry__2 
       (.CI(\I_4/multOp_carry__1_n_0 ),
        .CO({\I_4/multOp_carry__2_n_0 ,\I_4/multOp_carry__2_n_1 ,\I_4/multOp_carry__2_n_2 ,\I_4/multOp_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_4/plusOp_inferred__6_carry__1_n_5 }),
        .O({\I_4/multOp_carry__2_n_4 ,\I_4/multOp_carry__2_n_5 ,\I_4/multOp_carry__2_n_6 ,\I_4/multOp_carry__2_n_7 }),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,multOp_carry__2_i_1__0_n_0,multOp_carry__2_i_2__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_i_1 
       (.CI(\I_4/multOp_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[6] [10:8]}),
        .O({\I_4/multOp_i_1_n_4 ,\I_4/multOp_i_1_n_5 ,\I_4/multOp_i_1_n_6 ,\I_4/multOp_i_1_n_7 }),
        .S({\I_4/multOp_i_4_n_0 ,\I_4/multOp_i_5_n_0 ,\I_4/multOp_i_6_n_0 ,\I_4/multOp_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_10 
       (.I0(\sr_reg[6] [5]),
        .I1(\sr_reg[7] [5]),
        .O(\I_4/multOp_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_11 
       (.I0(\sr_reg[6] [4]),
        .I1(\sr_reg[7] [4]),
        .O(\I_4/multOp_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_12 
       (.I0(\sr_reg[6] [3]),
        .I1(\sr_reg[7] [3]),
        .O(\I_4/multOp_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_13 
       (.I0(\sr_reg[6] [2]),
        .I1(\sr_reg[7] [2]),
        .O(\I_4/multOp_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_14 
       (.I0(\sr_reg[6] [1]),
        .I1(\sr_reg[7] [1]),
        .O(\I_4/multOp_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_15 
       (.I0(\sr_reg[6] [0]),
        .I1(\sr_reg[7] [0]),
        .O(\I_4/multOp_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_i_2 
       (.CI(\I_4/multOp_i_3_n_0 ),
        .CO({\I_4/multOp_i_2_n_0 ,\I_4/multOp_i_2_n_1 ,\I_4/multOp_i_2_n_2 ,\I_4/multOp_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[6] [7:4]),
        .O({\I_4/multOp_i_2_n_4 ,\I_4/multOp_i_2_n_5 ,\I_4/multOp_i_2_n_6 ,\I_4/multOp_i_2_n_7 }),
        .S({\I_4/multOp_i_8_n_0 ,\I_4/multOp_i_9_n_0 ,\I_4/multOp_i_10_n_0 ,\I_4/multOp_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/multOp_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/multOp_i_3_n_0 ,\I_4/multOp_i_3_n_1 ,\I_4/multOp_i_3_n_2 ,\I_4/multOp_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[6] [3:0]),
        .O({\I_4/multOp_i_3_n_4 ,\I_4/multOp_i_3_n_5 ,\I_4/multOp_i_3_n_6 ,\I_4/multOp_i_3_n_7 }),
        .S({\I_4/multOp_i_12_n_0 ,\I_4/multOp_i_13_n_0 ,\I_4/multOp_i_14_n_0 ,\I_4/multOp_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_4 
       (.I0(\sr_reg[6] [11]),
        .I1(\sr_reg[7] [11]),
        .O(\I_4/multOp_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_5 
       (.I0(\sr_reg[6] [10]),
        .I1(\sr_reg[7] [10]),
        .O(\I_4/multOp_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_6 
       (.I0(\sr_reg[6] [9]),
        .I1(\sr_reg[7] [9]),
        .O(\I_4/multOp_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_7 
       (.I0(\sr_reg[6] [8]),
        .I1(\sr_reg[7] [8]),
        .O(\I_4/multOp_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_8 
       (.I0(\sr_reg[6] [7]),
        .I1(\sr_reg[7] [7]),
        .O(\I_4/multOp_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/multOp_i_9 
       (.I0(\sr_reg[6] [6]),
        .I1(\sr_reg[7] [6]),
        .O(\I_4/multOp_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\I_4/plusOp_inferred__7__62_carry__1_n_4 ),
        .Q(\I_4/output_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__4_n_6 ),
        .Q(\I_4/output_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__4_n_5 ),
        .Q(\I_4/output_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__2_n_7 ),
        .Q(\I_4/output_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__2_n_6 ),
        .Q(\I_4/output_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__2_n_5 ),
        .Q(\I_4/output_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__2_n_4 ),
        .Q(\I_4/output_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__3_n_7 ),
        .Q(\I_4/output_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__3_n_6 ),
        .Q(\I_4/output_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__3_n_5 ),
        .Q(\I_4/output_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__3_n_4 ),
        .Q(\I_4/output_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/output_reg[9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_4/plusOp_inferred__7__62_carry__4_n_7 ),
        .Q(\I_4/output_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/plusOp 
       (.A({\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_5 ,\I_4/plusOp_inferred__3_carry__1_n_6 ,\I_4/plusOp_inferred__3_carry__1_n_7 ,\I_4/plusOp_inferred__3_carry__0_n_4 ,\I_4/plusOp_inferred__3_carry__0_n_5 ,\I_4/plusOp_inferred__3_carry__0_n_6 ,\I_4/plusOp_inferred__3_carry__0_n_7 ,\I_4/plusOp_inferred__3_carry_n_4 ,\I_4/plusOp_inferred__3_carry_n_5 ,\I_4/plusOp_inferred__3_carry_n_6 ,\I_4/plusOp_inferred__3_carry_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_4/multOp_n_106 ,\I_4/multOp_n_107 ,\I_4/multOp_n_108 ,\I_4/multOp_n_109 ,\I_4/multOp_n_110 ,\I_4/multOp_n_111 ,\I_4/multOp_n_112 ,\I_4/multOp_n_113 ,\I_4/multOp_n_114 ,\I_4/multOp_n_115 ,\I_4/multOp_n_116 ,\I_4/multOp_n_117 ,\I_4/multOp_n_118 ,\I_4/multOp_n_119 ,\I_4/multOp_n_120 ,\I_4/multOp_n_121 ,\I_4/multOp_n_122 ,\I_4/multOp_n_123 ,\I_4/multOp_n_124 ,\I_4/multOp_n_125 ,\I_4/multOp_n_126 ,\I_4/multOp_n_127 ,\I_4/multOp_n_128 ,\I_4/multOp_n_129 ,\I_4/multOp_n_130 ,\I_4/multOp_n_131 ,\I_4/multOp_n_132 ,\I_4/multOp_n_133 ,\I_4/multOp_n_134 ,\I_4/multOp_n_135 ,\I_4/multOp_n_136 ,\I_4/multOp_n_137 ,\I_4/multOp_n_138 ,\I_4/multOp_n_139 ,\I_4/multOp_n_140 ,\I_4/multOp_n_141 ,\I_4/multOp_n_142 ,\I_4/multOp_n_143 ,\I_4/multOp_n_144 ,\I_4/multOp_n_145 ,\I_4/multOp_n_146 ,\I_4/multOp_n_147 ,\I_4/multOp_n_148 ,\I_4/multOp_n_149 ,\I_4/multOp_n_150 ,\I_4/multOp_n_151 ,\I_4/multOp_n_152 ,\I_4/multOp_n_153 }),
        .PCOUT({\I_4/plusOp_n_106 ,\I_4/plusOp_n_107 ,\I_4/plusOp_n_108 ,\I_4/plusOp_n_109 ,\I_4/plusOp_n_110 ,\I_4/plusOp_n_111 ,\I_4/plusOp_n_112 ,\I_4/plusOp_n_113 ,\I_4/plusOp_n_114 ,\I_4/plusOp_n_115 ,\I_4/plusOp_n_116 ,\I_4/plusOp_n_117 ,\I_4/plusOp_n_118 ,\I_4/plusOp_n_119 ,\I_4/plusOp_n_120 ,\I_4/plusOp_n_121 ,\I_4/plusOp_n_122 ,\I_4/plusOp_n_123 ,\I_4/plusOp_n_124 ,\I_4/plusOp_n_125 ,\I_4/plusOp_n_126 ,\I_4/plusOp_n_127 ,\I_4/plusOp_n_128 ,\I_4/plusOp_n_129 ,\I_4/plusOp_n_130 ,\I_4/plusOp_n_131 ,\I_4/plusOp_n_132 ,\I_4/plusOp_n_133 ,\I_4/plusOp_n_134 ,\I_4/plusOp_n_135 ,\I_4/plusOp_n_136 ,\I_4/plusOp_n_137 ,\I_4/plusOp_n_138 ,\I_4/plusOp_n_139 ,\I_4/plusOp_n_140 ,\I_4/plusOp_n_141 ,\I_4/plusOp_n_142 ,\I_4/plusOp_n_143 ,\I_4/plusOp_n_144 ,\I_4/plusOp_n_145 ,\I_4/plusOp_n_146 ,\I_4/plusOp_n_147 ,\I_4/plusOp_n_148 ,\I_4/plusOp_n_149 ,\I_4/plusOp_n_150 ,\I_4/plusOp_n_151 ,\I_4/plusOp_n_152 ,\I_4/plusOp_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/plusOp__0 
       (.A({\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_5 ,\I_4/plusOp__0_i_1_n_6 ,\I_4/plusOp__0_i_1_n_7 ,\I_4/plusOp__0_i_2_n_4 ,\I_4/plusOp__0_i_2_n_5 ,\I_4/plusOp__0_i_2_n_6 ,\I_4/plusOp__0_i_2_n_7 ,\I_4/plusOp__0_i_3_n_4 ,\I_4/plusOp__0_i_3_n_5 ,\I_4/plusOp__0_i_3_n_6 ,\I_4/plusOp__0_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_4/plusOp_n_106 ,\I_4/plusOp_n_107 ,\I_4/plusOp_n_108 ,\I_4/plusOp_n_109 ,\I_4/plusOp_n_110 ,\I_4/plusOp_n_111 ,\I_4/plusOp_n_112 ,\I_4/plusOp_n_113 ,\I_4/plusOp_n_114 ,\I_4/plusOp_n_115 ,\I_4/plusOp_n_116 ,\I_4/plusOp_n_117 ,\I_4/plusOp_n_118 ,\I_4/plusOp_n_119 ,\I_4/plusOp_n_120 ,\I_4/plusOp_n_121 ,\I_4/plusOp_n_122 ,\I_4/plusOp_n_123 ,\I_4/plusOp_n_124 ,\I_4/plusOp_n_125 ,\I_4/plusOp_n_126 ,\I_4/plusOp_n_127 ,\I_4/plusOp_n_128 ,\I_4/plusOp_n_129 ,\I_4/plusOp_n_130 ,\I_4/plusOp_n_131 ,\I_4/plusOp_n_132 ,\I_4/plusOp_n_133 ,\I_4/plusOp_n_134 ,\I_4/plusOp_n_135 ,\I_4/plusOp_n_136 ,\I_4/plusOp_n_137 ,\I_4/plusOp_n_138 ,\I_4/plusOp_n_139 ,\I_4/plusOp_n_140 ,\I_4/plusOp_n_141 ,\I_4/plusOp_n_142 ,\I_4/plusOp_n_143 ,\I_4/plusOp_n_144 ,\I_4/plusOp_n_145 ,\I_4/plusOp_n_146 ,\I_4/plusOp_n_147 ,\I_4/plusOp_n_148 ,\I_4/plusOp_n_149 ,\I_4/plusOp_n_150 ,\I_4/plusOp_n_151 ,\I_4/plusOp_n_152 ,\I_4/plusOp_n_153 }),
        .PCOUT({\I_4/plusOp__0_n_106 ,\I_4/plusOp__0_n_107 ,\I_4/plusOp__0_n_108 ,\I_4/plusOp__0_n_109 ,\I_4/plusOp__0_n_110 ,\I_4/plusOp__0_n_111 ,\I_4/plusOp__0_n_112 ,\I_4/plusOp__0_n_113 ,\I_4/plusOp__0_n_114 ,\I_4/plusOp__0_n_115 ,\I_4/plusOp__0_n_116 ,\I_4/plusOp__0_n_117 ,\I_4/plusOp__0_n_118 ,\I_4/plusOp__0_n_119 ,\I_4/plusOp__0_n_120 ,\I_4/plusOp__0_n_121 ,\I_4/plusOp__0_n_122 ,\I_4/plusOp__0_n_123 ,\I_4/plusOp__0_n_124 ,\I_4/plusOp__0_n_125 ,\I_4/plusOp__0_n_126 ,\I_4/plusOp__0_n_127 ,\I_4/plusOp__0_n_128 ,\I_4/plusOp__0_n_129 ,\I_4/plusOp__0_n_130 ,\I_4/plusOp__0_n_131 ,\I_4/plusOp__0_n_132 ,\I_4/plusOp__0_n_133 ,\I_4/plusOp__0_n_134 ,\I_4/plusOp__0_n_135 ,\I_4/plusOp__0_n_136 ,\I_4/plusOp__0_n_137 ,\I_4/plusOp__0_n_138 ,\I_4/plusOp__0_n_139 ,\I_4/plusOp__0_n_140 ,\I_4/plusOp__0_n_141 ,\I_4/plusOp__0_n_142 ,\I_4/plusOp__0_n_143 ,\I_4/plusOp__0_n_144 ,\I_4/plusOp__0_n_145 ,\I_4/plusOp__0_n_146 ,\I_4/plusOp__0_n_147 ,\I_4/plusOp__0_n_148 ,\I_4/plusOp__0_n_149 ,\I_4/plusOp__0_n_150 ,\I_4/plusOp__0_n_151 ,\I_4/plusOp__0_n_152 ,\I_4/plusOp__0_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__0_i_1 
       (.CI(\I_4/plusOp__0_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[5] [10:8]}),
        .O({\I_4/plusOp__0_i_1_n_4 ,\I_4/plusOp__0_i_1_n_5 ,\I_4/plusOp__0_i_1_n_6 ,\I_4/plusOp__0_i_1_n_7 }),
        .S({\I_4/plusOp__0_i_4_n_0 ,\I_4/plusOp__0_i_5_n_0 ,\I_4/plusOp__0_i_6_n_0 ,\I_4/plusOp__0_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_10 
       (.I0(\sr_reg[5] [5]),
        .I1(\sr_reg[8] [5]),
        .O(\I_4/plusOp__0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_11 
       (.I0(\sr_reg[5] [4]),
        .I1(\sr_reg[8] [4]),
        .O(\I_4/plusOp__0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_12 
       (.I0(\sr_reg[5] [3]),
        .I1(\sr_reg[8] [3]),
        .O(\I_4/plusOp__0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_13 
       (.I0(\sr_reg[5] [2]),
        .I1(\sr_reg[8] [2]),
        .O(\I_4/plusOp__0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_14 
       (.I0(\sr_reg[5] [1]),
        .I1(\sr_reg[8] [1]),
        .O(\I_4/plusOp__0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_15 
       (.I0(\sr_reg[5] [0]),
        .I1(\sr_reg[8] [0]),
        .O(\I_4/plusOp__0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__0_i_2 
       (.CI(\I_4/plusOp__0_i_3_n_0 ),
        .CO({\I_4/plusOp__0_i_2_n_0 ,\I_4/plusOp__0_i_2_n_1 ,\I_4/plusOp__0_i_2_n_2 ,\I_4/plusOp__0_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[5] [7:4]),
        .O({\I_4/plusOp__0_i_2_n_4 ,\I_4/plusOp__0_i_2_n_5 ,\I_4/plusOp__0_i_2_n_6 ,\I_4/plusOp__0_i_2_n_7 }),
        .S({\I_4/plusOp__0_i_8_n_0 ,\I_4/plusOp__0_i_9_n_0 ,\I_4/plusOp__0_i_10_n_0 ,\I_4/plusOp__0_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__0_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp__0_i_3_n_0 ,\I_4/plusOp__0_i_3_n_1 ,\I_4/plusOp__0_i_3_n_2 ,\I_4/plusOp__0_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[5] [3:0]),
        .O({\I_4/plusOp__0_i_3_n_4 ,\I_4/plusOp__0_i_3_n_5 ,\I_4/plusOp__0_i_3_n_6 ,\I_4/plusOp__0_i_3_n_7 }),
        .S({\I_4/plusOp__0_i_12_n_0 ,\I_4/plusOp__0_i_13_n_0 ,\I_4/plusOp__0_i_14_n_0 ,\I_4/plusOp__0_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_4 
       (.I0(\sr_reg[5] [11]),
        .I1(\sr_reg[8] [11]),
        .O(\I_4/plusOp__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_5 
       (.I0(\sr_reg[5] [10]),
        .I1(\sr_reg[8] [10]),
        .O(\I_4/plusOp__0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_6 
       (.I0(\sr_reg[5] [9]),
        .I1(\sr_reg[8] [9]),
        .O(\I_4/plusOp__0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_7 
       (.I0(\sr_reg[5] [8]),
        .I1(\sr_reg[8] [8]),
        .O(\I_4/plusOp__0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_8 
       (.I0(\sr_reg[5] [7]),
        .I1(\sr_reg[8] [7]),
        .O(\I_4/plusOp__0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__0_i_9 
       (.I0(\sr_reg[5] [6]),
        .I1(\sr_reg[8] [6]),
        .O(\I_4/plusOp__0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/plusOp__1 
       (.A({\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_5 ,\I_4/plusOp__1_i_1_n_6 ,\I_4/plusOp__1_i_1_n_7 ,\I_4/plusOp__1_i_2_n_4 ,\I_4/plusOp__1_i_2_n_5 ,\I_4/plusOp__1_i_2_n_6 ,\I_4/plusOp__1_i_2_n_7 ,\I_4/plusOp__1_i_3_n_4 ,\I_4/plusOp__1_i_3_n_5 ,\I_4/plusOp__1_i_3_n_6 ,\I_4/plusOp__1_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_4/plusOp__0_n_106 ,\I_4/plusOp__0_n_107 ,\I_4/plusOp__0_n_108 ,\I_4/plusOp__0_n_109 ,\I_4/plusOp__0_n_110 ,\I_4/plusOp__0_n_111 ,\I_4/plusOp__0_n_112 ,\I_4/plusOp__0_n_113 ,\I_4/plusOp__0_n_114 ,\I_4/plusOp__0_n_115 ,\I_4/plusOp__0_n_116 ,\I_4/plusOp__0_n_117 ,\I_4/plusOp__0_n_118 ,\I_4/plusOp__0_n_119 ,\I_4/plusOp__0_n_120 ,\I_4/plusOp__0_n_121 ,\I_4/plusOp__0_n_122 ,\I_4/plusOp__0_n_123 ,\I_4/plusOp__0_n_124 ,\I_4/plusOp__0_n_125 ,\I_4/plusOp__0_n_126 ,\I_4/plusOp__0_n_127 ,\I_4/plusOp__0_n_128 ,\I_4/plusOp__0_n_129 ,\I_4/plusOp__0_n_130 ,\I_4/plusOp__0_n_131 ,\I_4/plusOp__0_n_132 ,\I_4/plusOp__0_n_133 ,\I_4/plusOp__0_n_134 ,\I_4/plusOp__0_n_135 ,\I_4/plusOp__0_n_136 ,\I_4/plusOp__0_n_137 ,\I_4/plusOp__0_n_138 ,\I_4/plusOp__0_n_139 ,\I_4/plusOp__0_n_140 ,\I_4/plusOp__0_n_141 ,\I_4/plusOp__0_n_142 ,\I_4/plusOp__0_n_143 ,\I_4/plusOp__0_n_144 ,\I_4/plusOp__0_n_145 ,\I_4/plusOp__0_n_146 ,\I_4/plusOp__0_n_147 ,\I_4/plusOp__0_n_148 ,\I_4/plusOp__0_n_149 ,\I_4/plusOp__0_n_150 ,\I_4/plusOp__0_n_151 ,\I_4/plusOp__0_n_152 ,\I_4/plusOp__0_n_153 }),
        .PCOUT({\I_4/plusOp__1_n_106 ,\I_4/plusOp__1_n_107 ,\I_4/plusOp__1_n_108 ,\I_4/plusOp__1_n_109 ,\I_4/plusOp__1_n_110 ,\I_4/plusOp__1_n_111 ,\I_4/plusOp__1_n_112 ,\I_4/plusOp__1_n_113 ,\I_4/plusOp__1_n_114 ,\I_4/plusOp__1_n_115 ,\I_4/plusOp__1_n_116 ,\I_4/plusOp__1_n_117 ,\I_4/plusOp__1_n_118 ,\I_4/plusOp__1_n_119 ,\I_4/plusOp__1_n_120 ,\I_4/plusOp__1_n_121 ,\I_4/plusOp__1_n_122 ,\I_4/plusOp__1_n_123 ,\I_4/plusOp__1_n_124 ,\I_4/plusOp__1_n_125 ,\I_4/plusOp__1_n_126 ,\I_4/plusOp__1_n_127 ,\I_4/plusOp__1_n_128 ,\I_4/plusOp__1_n_129 ,\I_4/plusOp__1_n_130 ,\I_4/plusOp__1_n_131 ,\I_4/plusOp__1_n_132 ,\I_4/plusOp__1_n_133 ,\I_4/plusOp__1_n_134 ,\I_4/plusOp__1_n_135 ,\I_4/plusOp__1_n_136 ,\I_4/plusOp__1_n_137 ,\I_4/plusOp__1_n_138 ,\I_4/plusOp__1_n_139 ,\I_4/plusOp__1_n_140 ,\I_4/plusOp__1_n_141 ,\I_4/plusOp__1_n_142 ,\I_4/plusOp__1_n_143 ,\I_4/plusOp__1_n_144 ,\I_4/plusOp__1_n_145 ,\I_4/plusOp__1_n_146 ,\I_4/plusOp__1_n_147 ,\I_4/plusOp__1_n_148 ,\I_4/plusOp__1_n_149 ,\I_4/plusOp__1_n_150 ,\I_4/plusOp__1_n_151 ,\I_4/plusOp__1_n_152 ,\I_4/plusOp__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__1_i_1 
       (.CI(\I_4/plusOp__1_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[4] [10:8]}),
        .O({\I_4/plusOp__1_i_1_n_4 ,\I_4/plusOp__1_i_1_n_5 ,\I_4/plusOp__1_i_1_n_6 ,\I_4/plusOp__1_i_1_n_7 }),
        .S({\I_4/plusOp__1_i_4_n_0 ,\I_4/plusOp__1_i_5_n_0 ,\I_4/plusOp__1_i_6_n_0 ,\I_4/plusOp__1_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_10 
       (.I0(\sr_reg[4] [5]),
        .I1(\sr_reg[9] [5]),
        .O(\I_4/plusOp__1_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_11 
       (.I0(\sr_reg[4] [4]),
        .I1(\sr_reg[9] [4]),
        .O(\I_4/plusOp__1_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_12 
       (.I0(\sr_reg[4] [3]),
        .I1(\sr_reg[9] [3]),
        .O(\I_4/plusOp__1_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_13 
       (.I0(\sr_reg[4] [2]),
        .I1(\sr_reg[9] [2]),
        .O(\I_4/plusOp__1_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_14 
       (.I0(\sr_reg[4] [1]),
        .I1(\sr_reg[9] [1]),
        .O(\I_4/plusOp__1_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_15 
       (.I0(\sr_reg[4] [0]),
        .I1(\sr_reg[9] [0]),
        .O(\I_4/plusOp__1_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__1_i_2 
       (.CI(\I_4/plusOp__1_i_3_n_0 ),
        .CO({\I_4/plusOp__1_i_2_n_0 ,\I_4/plusOp__1_i_2_n_1 ,\I_4/plusOp__1_i_2_n_2 ,\I_4/plusOp__1_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[4] [7:4]),
        .O({\I_4/plusOp__1_i_2_n_4 ,\I_4/plusOp__1_i_2_n_5 ,\I_4/plusOp__1_i_2_n_6 ,\I_4/plusOp__1_i_2_n_7 }),
        .S({\I_4/plusOp__1_i_8_n_0 ,\I_4/plusOp__1_i_9_n_0 ,\I_4/plusOp__1_i_10_n_0 ,\I_4/plusOp__1_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__1_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp__1_i_3_n_0 ,\I_4/plusOp__1_i_3_n_1 ,\I_4/plusOp__1_i_3_n_2 ,\I_4/plusOp__1_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[4] [3:0]),
        .O({\I_4/plusOp__1_i_3_n_4 ,\I_4/plusOp__1_i_3_n_5 ,\I_4/plusOp__1_i_3_n_6 ,\I_4/plusOp__1_i_3_n_7 }),
        .S({\I_4/plusOp__1_i_12_n_0 ,\I_4/plusOp__1_i_13_n_0 ,\I_4/plusOp__1_i_14_n_0 ,\I_4/plusOp__1_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_4 
       (.I0(\sr_reg[4] [11]),
        .I1(\sr_reg[9] [11]),
        .O(\I_4/plusOp__1_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_5 
       (.I0(\sr_reg[4] [10]),
        .I1(\sr_reg[9] [10]),
        .O(\I_4/plusOp__1_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_6 
       (.I0(\sr_reg[4] [9]),
        .I1(\sr_reg[9] [9]),
        .O(\I_4/plusOp__1_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_7 
       (.I0(\sr_reg[4] [8]),
        .I1(\sr_reg[9] [8]),
        .O(\I_4/plusOp__1_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_8 
       (.I0(\sr_reg[4] [7]),
        .I1(\sr_reg[9] [7]),
        .O(\I_4/plusOp__1_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__1_i_9 
       (.I0(\sr_reg[4] [6]),
        .I1(\sr_reg[9] [6]),
        .O(\I_4/plusOp__1_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/plusOp__2 
       (.A({\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_5 ,\I_4/plusOp__2_i_1_n_6 ,\I_4/plusOp__2_i_1_n_7 ,\I_4/plusOp__2_i_2_n_4 ,\I_4/plusOp__2_i_2_n_5 ,\I_4/plusOp__2_i_2_n_6 ,\I_4/plusOp__2_i_2_n_7 ,\I_4/plusOp__2_i_3_n_4 ,\I_4/plusOp__2_i_3_n_5 ,\I_4/plusOp__2_i_3_n_6 ,\I_4/plusOp__2_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_4/plusOp__1_n_106 ,\I_4/plusOp__1_n_107 ,\I_4/plusOp__1_n_108 ,\I_4/plusOp__1_n_109 ,\I_4/plusOp__1_n_110 ,\I_4/plusOp__1_n_111 ,\I_4/plusOp__1_n_112 ,\I_4/plusOp__1_n_113 ,\I_4/plusOp__1_n_114 ,\I_4/plusOp__1_n_115 ,\I_4/plusOp__1_n_116 ,\I_4/plusOp__1_n_117 ,\I_4/plusOp__1_n_118 ,\I_4/plusOp__1_n_119 ,\I_4/plusOp__1_n_120 ,\I_4/plusOp__1_n_121 ,\I_4/plusOp__1_n_122 ,\I_4/plusOp__1_n_123 ,\I_4/plusOp__1_n_124 ,\I_4/plusOp__1_n_125 ,\I_4/plusOp__1_n_126 ,\I_4/plusOp__1_n_127 ,\I_4/plusOp__1_n_128 ,\I_4/plusOp__1_n_129 ,\I_4/plusOp__1_n_130 ,\I_4/plusOp__1_n_131 ,\I_4/plusOp__1_n_132 ,\I_4/plusOp__1_n_133 ,\I_4/plusOp__1_n_134 ,\I_4/plusOp__1_n_135 ,\I_4/plusOp__1_n_136 ,\I_4/plusOp__1_n_137 ,\I_4/plusOp__1_n_138 ,\I_4/plusOp__1_n_139 ,\I_4/plusOp__1_n_140 ,\I_4/plusOp__1_n_141 ,\I_4/plusOp__1_n_142 ,\I_4/plusOp__1_n_143 ,\I_4/plusOp__1_n_144 ,\I_4/plusOp__1_n_145 ,\I_4/plusOp__1_n_146 ,\I_4/plusOp__1_n_147 ,\I_4/plusOp__1_n_148 ,\I_4/plusOp__1_n_149 ,\I_4/plusOp__1_n_150 ,\I_4/plusOp__1_n_151 ,\I_4/plusOp__1_n_152 ,\I_4/plusOp__1_n_153 }),
        .PCOUT({\I_4/plusOp__2_n_106 ,\I_4/plusOp__2_n_107 ,\I_4/plusOp__2_n_108 ,\I_4/plusOp__2_n_109 ,\I_4/plusOp__2_n_110 ,\I_4/plusOp__2_n_111 ,\I_4/plusOp__2_n_112 ,\I_4/plusOp__2_n_113 ,\I_4/plusOp__2_n_114 ,\I_4/plusOp__2_n_115 ,\I_4/plusOp__2_n_116 ,\I_4/plusOp__2_n_117 ,\I_4/plusOp__2_n_118 ,\I_4/plusOp__2_n_119 ,\I_4/plusOp__2_n_120 ,\I_4/plusOp__2_n_121 ,\I_4/plusOp__2_n_122 ,\I_4/plusOp__2_n_123 ,\I_4/plusOp__2_n_124 ,\I_4/plusOp__2_n_125 ,\I_4/plusOp__2_n_126 ,\I_4/plusOp__2_n_127 ,\I_4/plusOp__2_n_128 ,\I_4/plusOp__2_n_129 ,\I_4/plusOp__2_n_130 ,\I_4/plusOp__2_n_131 ,\I_4/plusOp__2_n_132 ,\I_4/plusOp__2_n_133 ,\I_4/plusOp__2_n_134 ,\I_4/plusOp__2_n_135 ,\I_4/plusOp__2_n_136 ,\I_4/plusOp__2_n_137 ,\I_4/plusOp__2_n_138 ,\I_4/plusOp__2_n_139 ,\I_4/plusOp__2_n_140 ,\I_4/plusOp__2_n_141 ,\I_4/plusOp__2_n_142 ,\I_4/plusOp__2_n_143 ,\I_4/plusOp__2_n_144 ,\I_4/plusOp__2_n_145 ,\I_4/plusOp__2_n_146 ,\I_4/plusOp__2_n_147 ,\I_4/plusOp__2_n_148 ,\I_4/plusOp__2_n_149 ,\I_4/plusOp__2_n_150 ,\I_4/plusOp__2_n_151 ,\I_4/plusOp__2_n_152 ,\I_4/plusOp__2_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__2_i_1 
       (.CI(\I_4/plusOp__2_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[3] [10:8]}),
        .O({\I_4/plusOp__2_i_1_n_4 ,\I_4/plusOp__2_i_1_n_5 ,\I_4/plusOp__2_i_1_n_6 ,\I_4/plusOp__2_i_1_n_7 }),
        .S({\I_4/plusOp__2_i_4_n_0 ,\I_4/plusOp__2_i_5_n_0 ,\I_4/plusOp__2_i_6_n_0 ,\I_4/plusOp__2_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_10 
       (.I0(\sr_reg[3] [5]),
        .I1(\sr_reg[10] [5]),
        .O(\I_4/plusOp__2_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_11 
       (.I0(\sr_reg[3] [4]),
        .I1(\sr_reg[10] [4]),
        .O(\I_4/plusOp__2_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_12 
       (.I0(\sr_reg[3] [3]),
        .I1(\sr_reg[10] [3]),
        .O(\I_4/plusOp__2_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_13 
       (.I0(\sr_reg[3] [2]),
        .I1(\sr_reg[10] [2]),
        .O(\I_4/plusOp__2_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_14 
       (.I0(\sr_reg[3] [1]),
        .I1(\sr_reg[10] [1]),
        .O(\I_4/plusOp__2_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_15 
       (.I0(\sr_reg[3] [0]),
        .I1(\sr_reg[10] [0]),
        .O(\I_4/plusOp__2_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__2_i_2 
       (.CI(\I_4/plusOp__2_i_3_n_0 ),
        .CO({\I_4/plusOp__2_i_2_n_0 ,\I_4/plusOp__2_i_2_n_1 ,\I_4/plusOp__2_i_2_n_2 ,\I_4/plusOp__2_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[3] [7:4]),
        .O({\I_4/plusOp__2_i_2_n_4 ,\I_4/plusOp__2_i_2_n_5 ,\I_4/plusOp__2_i_2_n_6 ,\I_4/plusOp__2_i_2_n_7 }),
        .S({\I_4/plusOp__2_i_8_n_0 ,\I_4/plusOp__2_i_9_n_0 ,\I_4/plusOp__2_i_10_n_0 ,\I_4/plusOp__2_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__2_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp__2_i_3_n_0 ,\I_4/plusOp__2_i_3_n_1 ,\I_4/plusOp__2_i_3_n_2 ,\I_4/plusOp__2_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[3] [3:0]),
        .O({\I_4/plusOp__2_i_3_n_4 ,\I_4/plusOp__2_i_3_n_5 ,\I_4/plusOp__2_i_3_n_6 ,\I_4/plusOp__2_i_3_n_7 }),
        .S({\I_4/plusOp__2_i_12_n_0 ,\I_4/plusOp__2_i_13_n_0 ,\I_4/plusOp__2_i_14_n_0 ,\I_4/plusOp__2_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_4 
       (.I0(\sr_reg[3] [11]),
        .I1(\sr_reg[10] [11]),
        .O(\I_4/plusOp__2_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_5 
       (.I0(\sr_reg[3] [10]),
        .I1(\sr_reg[10] [10]),
        .O(\I_4/plusOp__2_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_6 
       (.I0(\sr_reg[3] [9]),
        .I1(\sr_reg[10] [9]),
        .O(\I_4/plusOp__2_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_7 
       (.I0(\sr_reg[3] [8]),
        .I1(\sr_reg[10] [8]),
        .O(\I_4/plusOp__2_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_8 
       (.I0(\sr_reg[3] [7]),
        .I1(\sr_reg[10] [7]),
        .O(\I_4/plusOp__2_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__2_i_9 
       (.I0(\sr_reg[3] [6]),
        .I1(\sr_reg[10] [6]),
        .O(\I_4/plusOp__2_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_4/plusOp__3 
       (.A({\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_5 ,\I_4/plusOp__3_i_1_n_6 ,\I_4/plusOp__3_i_1_n_7 ,\I_4/plusOp__3_i_2_n_4 ,\I_4/plusOp__3_i_2_n_5 ,\I_4/plusOp__3_i_2_n_6 ,\I_4/plusOp__3_i_2_n_7 ,\I_4/plusOp__3_i_3_n_4 ,\I_4/plusOp__3_i_3_n_5 ,\I_4/plusOp__3_i_3_n_6 ,\I_4/plusOp__3_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\I_4/plusOp__3_n_58 ,\I_4/plusOp__3_n_59 ,\I_4/plusOp__3_n_60 ,\I_4/plusOp__3_n_61 ,\I_4/plusOp__3_n_62 ,\I_4/plusOp__3_n_63 ,\I_4/plusOp__3_n_64 ,\I_4/plusOp__3_n_65 ,\I_4/plusOp__3_n_66 ,\I_4/plusOp__3_n_67 ,\I_4/plusOp__3_n_68 ,\I_4/plusOp__3_n_69 ,\I_4/plusOp__3_n_70 ,\I_4/plusOp__3_n_71 ,\I_4/plusOp__3_n_72 ,\I_4/plusOp__3_n_73 ,\I_4/plusOp__3_n_74 ,\I_4/plusOp__3_n_75 ,\I_4/plusOp__3_n_76 ,\I_4/plusOp__3_n_77 ,\I_4/plusOp__3_n_78 ,\I_4/plusOp__3_n_79 ,\I_4/plusOp__3_n_80 ,\I_4/plusOp__3_n_81 ,\I_4/plusOp__3_n_82 ,\I_4/plusOp__3_n_83 ,\I_4/plusOp__3_n_84 ,\I_4/plusOp__3_n_85 ,\I_4/plusOp__3_n_86 ,\I_4/plusOp__3_n_87 ,\I_4/plusOp__3_n_88 ,\I_4/plusOp__3_n_89 ,\I_4/plusOp__3_n_90 ,\I_4/plusOp__3_n_91 ,\I_4/plusOp__3_n_92 ,\I_4/plusOp__3_n_93 ,\I_4/plusOp__3_n_94 ,\I_4/plusOp__3_n_95 ,\I_4/plusOp__3_n_96 ,\I_4/plusOp__3_n_97 ,\I_4/plusOp__3_n_98 ,\I_4/plusOp__3_n_99 ,\I_4/plusOp__3_n_100 ,\I_4/plusOp__3_n_101 ,\I_4/plusOp__3_n_102 ,\I_4/plusOp__3_n_103 ,\I_4/plusOp__3_n_104 ,\I_4/plusOp__3_n_105 }),
        .PCIN({\I_4/plusOp__2_n_106 ,\I_4/plusOp__2_n_107 ,\I_4/plusOp__2_n_108 ,\I_4/plusOp__2_n_109 ,\I_4/plusOp__2_n_110 ,\I_4/plusOp__2_n_111 ,\I_4/plusOp__2_n_112 ,\I_4/plusOp__2_n_113 ,\I_4/plusOp__2_n_114 ,\I_4/plusOp__2_n_115 ,\I_4/plusOp__2_n_116 ,\I_4/plusOp__2_n_117 ,\I_4/plusOp__2_n_118 ,\I_4/plusOp__2_n_119 ,\I_4/plusOp__2_n_120 ,\I_4/plusOp__2_n_121 ,\I_4/plusOp__2_n_122 ,\I_4/plusOp__2_n_123 ,\I_4/plusOp__2_n_124 ,\I_4/plusOp__2_n_125 ,\I_4/plusOp__2_n_126 ,\I_4/plusOp__2_n_127 ,\I_4/plusOp__2_n_128 ,\I_4/plusOp__2_n_129 ,\I_4/plusOp__2_n_130 ,\I_4/plusOp__2_n_131 ,\I_4/plusOp__2_n_132 ,\I_4/plusOp__2_n_133 ,\I_4/plusOp__2_n_134 ,\I_4/plusOp__2_n_135 ,\I_4/plusOp__2_n_136 ,\I_4/plusOp__2_n_137 ,\I_4/plusOp__2_n_138 ,\I_4/plusOp__2_n_139 ,\I_4/plusOp__2_n_140 ,\I_4/plusOp__2_n_141 ,\I_4/plusOp__2_n_142 ,\I_4/plusOp__2_n_143 ,\I_4/plusOp__2_n_144 ,\I_4/plusOp__2_n_145 ,\I_4/plusOp__2_n_146 ,\I_4/plusOp__2_n_147 ,\I_4/plusOp__2_n_148 ,\I_4/plusOp__2_n_149 ,\I_4/plusOp__2_n_150 ,\I_4/plusOp__2_n_151 ,\I_4/plusOp__2_n_152 ,\I_4/plusOp__2_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__3_i_1 
       (.CI(\I_4/plusOp__3_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[2] [10:8]}),
        .O({\I_4/plusOp__3_i_1_n_4 ,\I_4/plusOp__3_i_1_n_5 ,\I_4/plusOp__3_i_1_n_6 ,\I_4/plusOp__3_i_1_n_7 }),
        .S({\I_4/plusOp__3_i_4_n_0 ,\I_4/plusOp__3_i_5_n_0 ,\I_4/plusOp__3_i_6_n_0 ,\I_4/plusOp__3_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_10 
       (.I0(\sr_reg[2] [5]),
        .I1(\sr_reg[11] [5]),
        .O(\I_4/plusOp__3_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_11 
       (.I0(\sr_reg[2] [4]),
        .I1(\sr_reg[11] [4]),
        .O(\I_4/plusOp__3_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_12 
       (.I0(\sr_reg[2] [3]),
        .I1(\sr_reg[11] [3]),
        .O(\I_4/plusOp__3_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_13 
       (.I0(\sr_reg[2] [2]),
        .I1(\sr_reg[11] [2]),
        .O(\I_4/plusOp__3_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_14 
       (.I0(\sr_reg[2] [1]),
        .I1(\sr_reg[11] [1]),
        .O(\I_4/plusOp__3_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_15 
       (.I0(\sr_reg[2] [0]),
        .I1(\sr_reg[11] [0]),
        .O(\I_4/plusOp__3_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__3_i_2 
       (.CI(\I_4/plusOp__3_i_3_n_0 ),
        .CO({\I_4/plusOp__3_i_2_n_0 ,\I_4/plusOp__3_i_2_n_1 ,\I_4/plusOp__3_i_2_n_2 ,\I_4/plusOp__3_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[2] [7:4]),
        .O({\I_4/plusOp__3_i_2_n_4 ,\I_4/plusOp__3_i_2_n_5 ,\I_4/plusOp__3_i_2_n_6 ,\I_4/plusOp__3_i_2_n_7 }),
        .S({\I_4/plusOp__3_i_8_n_0 ,\I_4/plusOp__3_i_9_n_0 ,\I_4/plusOp__3_i_10_n_0 ,\I_4/plusOp__3_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp__3_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp__3_i_3_n_0 ,\I_4/plusOp__3_i_3_n_1 ,\I_4/plusOp__3_i_3_n_2 ,\I_4/plusOp__3_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[2] [3:0]),
        .O({\I_4/plusOp__3_i_3_n_4 ,\I_4/plusOp__3_i_3_n_5 ,\I_4/plusOp__3_i_3_n_6 ,\I_4/plusOp__3_i_3_n_7 }),
        .S({\I_4/plusOp__3_i_12_n_0 ,\I_4/plusOp__3_i_13_n_0 ,\I_4/plusOp__3_i_14_n_0 ,\I_4/plusOp__3_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_4 
       (.I0(\sr_reg[2] [11]),
        .I1(\sr_reg[11] [11]),
        .O(\I_4/plusOp__3_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_5 
       (.I0(\sr_reg[2] [10]),
        .I1(\sr_reg[11] [10]),
        .O(\I_4/plusOp__3_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_6 
       (.I0(\sr_reg[2] [9]),
        .I1(\sr_reg[11] [9]),
        .O(\I_4/plusOp__3_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_7 
       (.I0(\sr_reg[2] [8]),
        .I1(\sr_reg[11] [8]),
        .O(\I_4/plusOp__3_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_8 
       (.I0(\sr_reg[2] [7]),
        .I1(\sr_reg[11] [7]),
        .O(\I_4/plusOp__3_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_4/plusOp__3_i_9 
       (.I0(\sr_reg[2] [6]),
        .I1(\sr_reg[11] [6]),
        .O(\I_4/plusOp__3_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__3_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp_inferred__3_carry_n_0 ,\I_4/plusOp_inferred__3_carry_n_1 ,\I_4/plusOp_inferred__3_carry_n_2 ,\I_4/plusOp_inferred__3_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[14] [3:0]),
        .O({\I_4/plusOp_inferred__3_carry_n_4 ,\I_4/plusOp_inferred__3_carry_n_5 ,\I_4/plusOp_inferred__3_carry_n_6 ,\I_4/plusOp_inferred__3_carry_n_7 }),
        .S({plusOp_inferred__3_carry_i_1__0_n_0,plusOp_inferred__3_carry_i_2__0_n_0,plusOp_inferred__3_carry_i_3__0_n_0,plusOp_inferred__3_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__3_carry__0 
       (.CI(\I_4/plusOp_inferred__3_carry_n_0 ),
        .CO({\I_4/plusOp_inferred__3_carry__0_n_0 ,\I_4/plusOp_inferred__3_carry__0_n_1 ,\I_4/plusOp_inferred__3_carry__0_n_2 ,\I_4/plusOp_inferred__3_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[14] [7:4]),
        .O({\I_4/plusOp_inferred__3_carry__0_n_4 ,\I_4/plusOp_inferred__3_carry__0_n_5 ,\I_4/plusOp_inferred__3_carry__0_n_6 ,\I_4/plusOp_inferred__3_carry__0_n_7 }),
        .S({plusOp_inferred__3_carry__0_i_1__0_n_0,plusOp_inferred__3_carry__0_i_2__0_n_0,plusOp_inferred__3_carry__0_i_3__0_n_0,plusOp_inferred__3_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__3_carry__1 
       (.CI(\I_4/plusOp_inferred__3_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[14] [10:8]}),
        .O({\I_4/plusOp_inferred__3_carry__1_n_4 ,\I_4/plusOp_inferred__3_carry__1_n_5 ,\I_4/plusOp_inferred__3_carry__1_n_6 ,\I_4/plusOp_inferred__3_carry__1_n_7 }),
        .S({plusOp_inferred__3_carry__1_i_1__0_n_0,plusOp_inferred__3_carry__1_i_2__0_n_0,plusOp_inferred__3_carry__1_i_3__0_n_0,plusOp_inferred__3_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__5_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp_inferred__5_carry_n_0 ,\I_4/plusOp_inferred__5_carry_n_1 ,\I_4/plusOp_inferred__5_carry_n_2 ,\I_4/plusOp_inferred__5_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[1] [3:0]),
        .O(\I_4/multOp__0 [3:0]),
        .S({plusOp_inferred__5_carry_i_1__0_n_0,plusOp_inferred__5_carry_i_2__0_n_0,plusOp_inferred__5_carry_i_3__0_n_0,plusOp_inferred__5_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__5_carry__0 
       (.CI(\I_4/plusOp_inferred__5_carry_n_0 ),
        .CO({\I_4/plusOp_inferred__5_carry__0_n_0 ,\I_4/plusOp_inferred__5_carry__0_n_1 ,\I_4/plusOp_inferred__5_carry__0_n_2 ,\I_4/plusOp_inferred__5_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[1] [7:4]),
        .O(\I_4/multOp__0 [7:4]),
        .S({plusOp_inferred__5_carry__0_i_1__0_n_0,plusOp_inferred__5_carry__0_i_2__0_n_0,plusOp_inferred__5_carry__0_i_3__0_n_0,plusOp_inferred__5_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__5_carry__1 
       (.CI(\I_4/plusOp_inferred__5_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[1] [10:8]}),
        .O(\I_4/multOp__0 [11:8]),
        .S({plusOp_inferred__5_carry__1_i_1__0_n_0,plusOp_inferred__5_carry__1_i_2__0_n_0,plusOp_inferred__5_carry__1_i_3__0_n_0,plusOp_inferred__5_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__6_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp_inferred__6_carry_n_0 ,\I_4/plusOp_inferred__6_carry_n_1 ,\I_4/plusOp_inferred__6_carry_n_2 ,\I_4/plusOp_inferred__6_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[0] [3:0]),
        .O({\I_4/plusOp_inferred__6_carry_n_4 ,\I_4/plusOp_inferred__6_carry_n_5 ,\I_4/plusOp_inferred__6_carry_n_6 ,\I_4/plusOp_inferred__6_carry_n_7 }),
        .S({plusOp_inferred__6_carry_i_1__0_n_0,plusOp_inferred__6_carry_i_2__0_n_0,plusOp_inferred__6_carry_i_3__0_n_0,plusOp_inferred__6_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__6_carry__0 
       (.CI(\I_4/plusOp_inferred__6_carry_n_0 ),
        .CO({\I_4/plusOp_inferred__6_carry__0_n_0 ,\I_4/plusOp_inferred__6_carry__0_n_1 ,\I_4/plusOp_inferred__6_carry__0_n_2 ,\I_4/plusOp_inferred__6_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\sr_reg[0] [7:4]),
        .O({\I_4/plusOp_inferred__6_carry__0_n_4 ,\I_4/plusOp_inferred__6_carry__0_n_5 ,\I_4/plusOp_inferred__6_carry__0_n_6 ,\I_4/plusOp_inferred__6_carry__0_n_7 }),
        .S({plusOp_inferred__6_carry__0_i_1__0_n_0,plusOp_inferred__6_carry__0_i_2__0_n_0,plusOp_inferred__6_carry__0_i_3__0_n_0,plusOp_inferred__6_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__6_carry__1 
       (.CI(\I_4/plusOp_inferred__6_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\sr_reg[0] [10:8]}),
        .O({\I_4/plusOp_inferred__6_carry__1_n_4 ,\I_4/plusOp_inferred__6_carry__1_n_5 ,\I_4/plusOp_inferred__6_carry__1_n_6 ,\I_4/plusOp_inferred__6_carry__1_n_7 }),
        .S({plusOp_inferred__6_carry__1_i_1__0_n_0,plusOp_inferred__6_carry__1_i_2__0_n_0,plusOp_inferred__6_carry__1_i_3__0_n_0,plusOp_inferred__6_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp_inferred__7__62_carry_n_0 ,\I_4/plusOp_inferred__7__62_carry_n_1 ,\I_4/plusOp_inferred__7__62_carry_n_2 ,\I_4/plusOp_inferred__7__62_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(multOp0[3:0]),
        .S({plusOp_inferred__7__62_carry_i_1__0_n_0,plusOp_inferred__7__62_carry_i_2__0_n_0,plusOp_inferred__7__62_carry_i_3__0_n_0,plusOp_inferred__7__62_carry_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry__0 
       (.CI(\I_4/plusOp_inferred__7__62_carry_n_0 ),
        .CO({\I_4/plusOp_inferred__7__62_carry__0_n_0 ,\I_4/plusOp_inferred__7__62_carry__0_n_1 ,\I_4/plusOp_inferred__7__62_carry__0_n_2 ,\I_4/plusOp_inferred__7__62_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(multOp0[7:4]),
        .S({plusOp_inferred__7__62_carry__0_i_1__0_n_0,plusOp_inferred__7__62_carry__0_i_2__0_n_0,plusOp_inferred__7__62_carry__0_i_3__0_n_0,plusOp_inferred__7__62_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry__1 
       (.CI(\I_4/plusOp_inferred__7__62_carry__0_n_0 ),
        .CO({\I_4/plusOp_inferred__7__62_carry__1_n_0 ,\I_4/plusOp_inferred__7__62_carry__1_n_1 ,\I_4/plusOp_inferred__7__62_carry__1_n_2 ,\I_4/plusOp_inferred__7__62_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(multOp0[11:8]),
        .O({\I_4/plusOp_inferred__7__62_carry__1_n_4 ,\I_4/plusOp_inferred__7__62_carry__1_n_5 ,\I_4/plusOp_inferred__7__62_carry__1_n_6 ,\I_4/plusOp_inferred__7__62_carry__1_n_7 }),
        .S({plusOp_inferred__7__62_carry__1_i_1__0_n_0,plusOp_inferred__7__62_carry__1_i_2__0_n_0,plusOp_inferred__7__62_carry__1_i_3__0_n_0,plusOp_inferred__7__62_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry__2 
       (.CI(\I_4/plusOp_inferred__7__62_carry__1_n_0 ),
        .CO({\I_4/plusOp_inferred__7__62_carry__2_n_0 ,\I_4/plusOp_inferred__7__62_carry__2_n_1 ,\I_4/plusOp_inferred__7__62_carry__2_n_2 ,\I_4/plusOp_inferred__7__62_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({plusOp_inferred__7__62_carry__2_i_1__0_n_0,multOp0[14:12]}),
        .O({\I_4/plusOp_inferred__7__62_carry__2_n_4 ,\I_4/plusOp_inferred__7__62_carry__2_n_5 ,\I_4/plusOp_inferred__7__62_carry__2_n_6 ,\I_4/plusOp_inferred__7__62_carry__2_n_7 }),
        .S({plusOp_inferred__7__62_carry__2_i_2__0_n_0,plusOp_inferred__7__62_carry__2_i_3__0_n_0,plusOp_inferred__7__62_carry__2_i_4__0_n_0,plusOp_inferred__7__62_carry__2_i_5__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry__3 
       (.CI(\I_4/plusOp_inferred__7__62_carry__2_n_0 ),
        .CO({\I_4/plusOp_inferred__7__62_carry__3_n_0 ,\I_4/plusOp_inferred__7__62_carry__3_n_1 ,\I_4/plusOp_inferred__7__62_carry__3_n_2 ,\I_4/plusOp_inferred__7__62_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(C__0[18:15]),
        .O({\I_4/plusOp_inferred__7__62_carry__3_n_4 ,\I_4/plusOp_inferred__7__62_carry__3_n_5 ,\I_4/plusOp_inferred__7__62_carry__3_n_6 ,\I_4/plusOp_inferred__7__62_carry__3_n_7 }),
        .S({plusOp_inferred__7__62_carry__3_i_1__0_n_0,plusOp_inferred__7__62_carry__3_i_2__0_n_0,plusOp_inferred__7__62_carry__3_i_3__0_n_0,plusOp_inferred__7__62_carry__3_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7__62_carry__4 
       (.CI(\I_4/plusOp_inferred__7__62_carry__3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,C__0[20:19]}),
        .O({\I_4/plusOp_inferred__7__62_carry__4_n_4 ,\I_4/plusOp_inferred__7__62_carry__4_n_5 ,\I_4/plusOp_inferred__7__62_carry__4_n_6 ,\I_4/plusOp_inferred__7__62_carry__4_n_7 }),
        .S({\<const0>__0__0 ,plusOp_inferred__7__62_carry__4_i_1__0_n_0,plusOp_inferred__7__62_carry__4_i_2__0_n_0,plusOp_inferred__7__62_carry__4_i_3__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_4/plusOp_inferred__7_carry_n_0 ,\I_4/plusOp_inferred__7_carry_n_1 ,\I_4/plusOp_inferred__7_carry_n_2 ,\I_4/plusOp_inferred__7_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/multOp__0 [2:0],\<const0>__0__0 }),
        .O(C__0[4:1]),
        .S({plusOp_inferred__7_carry_i_1__0_n_0,plusOp_inferred__7_carry_i_2__0_n_0,plusOp_inferred__7_carry_i_3__0_n_0,\I_4/plusOp__3_n_104 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry__0 
       (.CI(\I_4/plusOp_inferred__7_carry_n_0 ),
        .CO({\I_4/plusOp_inferred__7_carry__0_n_0 ,\I_4/plusOp_inferred__7_carry__0_n_1 ,\I_4/plusOp_inferred__7_carry__0_n_2 ,\I_4/plusOp_inferred__7_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_4/multOp__0 [6:3]),
        .O(C__0[8:5]),
        .S({plusOp_inferred__7_carry__0_i_1__0_n_0,plusOp_inferred__7_carry__0_i_2__0_n_0,plusOp_inferred__7_carry__0_i_3__0_n_0,plusOp_inferred__7_carry__0_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry__1 
       (.CI(\I_4/plusOp_inferred__7_carry__0_n_0 ),
        .CO({\I_4/plusOp_inferred__7_carry__1_n_0 ,\I_4/plusOp_inferred__7_carry__1_n_1 ,\I_4/plusOp_inferred__7_carry__1_n_2 ,\I_4/plusOp_inferred__7_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_4/multOp__0 [10:7]),
        .O(C__0[12:9]),
        .S({plusOp_inferred__7_carry__1_i_1__0_n_0,plusOp_inferred__7_carry__1_i_2__0_n_0,plusOp_inferred__7_carry__1_i_3__0_n_0,plusOp_inferred__7_carry__1_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry__2 
       (.CI(\I_4/plusOp_inferred__7_carry__1_n_0 ),
        .CO({\I_4/plusOp_inferred__7_carry__2_n_0 ,\I_4/plusOp_inferred__7_carry__2_n_1 ,\I_4/plusOp_inferred__7_carry__2_n_2 ,\I_4/plusOp_inferred__7_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/plusOp__3_n_90 ,\I_4/plusOp__3_n_91 ,\I_4/plusOp__3_n_92 ,plusOp_inferred__7_carry__2_i_1__0_n_0}),
        .O(C__0[16:13]),
        .S({plusOp_inferred__7_carry__2_i_2__0_n_0,plusOp_inferred__7_carry__2_i_3__0_n_0,plusOp_inferred__7_carry__2_i_4__0_n_0,plusOp_inferred__7_carry__2_i_5__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry__3 
       (.CI(\I_4/plusOp_inferred__7_carry__2_n_0 ),
        .CO({\I_4/plusOp_inferred__7_carry__3_n_0 ,\I_4/plusOp_inferred__7_carry__3_n_1 ,\I_4/plusOp_inferred__7_carry__3_n_2 ,\I_4/plusOp_inferred__7_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_4/plusOp__3_n_86 ,\I_4/plusOp__3_n_87 ,\I_4/plusOp__3_n_88 ,\I_4/plusOp__3_n_89 }),
        .O(C__0[20:17]),
        .S({plusOp_inferred__7_carry__3_i_1__0_n_0,plusOp_inferred__7_carry__3_i_2__0_n_0,plusOp_inferred__7_carry__3_i_3__0_n_0,plusOp_inferred__7_carry__3_i_4__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_4/plusOp_inferred__7_carry__4 
       (.CI(\I_4/plusOp_inferred__7_carry__3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_4/plusOp__3_n_85 }),
        .O({\I_4/plusOp_inferred__7_carry__4_n_4 ,\I_4/plusOp_inferred__7_carry__4_n_5 ,C__0[22:21]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,plusOp_inferred__7_carry__4_i_1__0_n_0,plusOp_inferred__7_carry__4_i_2__0_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [0]),
        .Q(\sr_reg[0] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [10]),
        .Q(\sr_reg[0] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [11]),
        .Q(\sr_reg[0] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [1]),
        .Q(\sr_reg[0] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [2]),
        .Q(\sr_reg[0] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [3]),
        .Q(\sr_reg[0] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [4]),
        .Q(\sr_reg[0] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [5]),
        .Q(\sr_reg[0] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [6]),
        .Q(\sr_reg[0] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [7]),
        .Q(\sr_reg[0] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [8]),
        .Q(\sr_reg[0] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[0][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\input [9]),
        .Q(\sr_reg[0] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [0]),
        .Q(\sr_reg[10] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [10]),
        .Q(\sr_reg[10] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [11]),
        .Q(\sr_reg[10] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [1]),
        .Q(\sr_reg[10] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [2]),
        .Q(\sr_reg[10] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [3]),
        .Q(\sr_reg[10] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[9] [4]),
        .Q(\sr_reg[10] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[9] [5]),
        .Q(\sr_reg[10] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[9] [6]),
        .Q(\sr_reg[10] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[9] [7]),
        .Q(\sr_reg[10] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [8]),
        .Q(\sr_reg[10] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[10][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[9] [9]),
        .Q(\sr_reg[10] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [0]),
        .Q(\sr_reg[11] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[10] [10]),
        .Q(\sr_reg[11] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[10] [11]),
        .Q(\sr_reg[11] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [1]),
        .Q(\sr_reg[11] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [2]),
        .Q(\sr_reg[11] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [3]),
        .Q(\sr_reg[11] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [4]),
        .Q(\sr_reg[11] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [5]),
        .Q(\sr_reg[11] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [6]),
        .Q(\sr_reg[11] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[10] [7]),
        .Q(\sr_reg[11] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[10] [8]),
        .Q(\sr_reg[11] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[11][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[10] [9]),
        .Q(\sr_reg[11] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [0]),
        .Q(\sr_reg[12] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [10]),
        .Q(\sr_reg[12] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [11]),
        .Q(\sr_reg[12] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [1]),
        .Q(\sr_reg[12] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [2]),
        .Q(\sr_reg[12] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [3]),
        .Q(\sr_reg[12] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [4]),
        .Q(\sr_reg[12] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [5]),
        .Q(\sr_reg[12] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [6]),
        .Q(\sr_reg[12] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [7]),
        .Q(\sr_reg[12] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [8]),
        .Q(\sr_reg[12] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[12][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[11] [9]),
        .Q(\sr_reg[12] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [0]),
        .Q(\sr_reg[13] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [10]),
        .Q(\sr_reg[13] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [11]),
        .Q(\sr_reg[13] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [1]),
        .Q(\sr_reg[13] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [2]),
        .Q(\sr_reg[13] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [3]),
        .Q(\sr_reg[13] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [4]),
        .Q(\sr_reg[13] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [5]),
        .Q(\sr_reg[13] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [6]),
        .Q(\sr_reg[13] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [7]),
        .Q(\sr_reg[13] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [8]),
        .Q(\sr_reg[13] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[13][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[12] [9]),
        .Q(\sr_reg[13] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [0]),
        .Q(\sr_reg[14] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [10]),
        .Q(\sr_reg[14] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [11]),
        .Q(\sr_reg[14] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [1]),
        .Q(\sr_reg[14] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [2]),
        .Q(\sr_reg[14] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [3]),
        .Q(\sr_reg[14] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [4]),
        .Q(\sr_reg[14] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [5]),
        .Q(\sr_reg[14] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [6]),
        .Q(\sr_reg[14] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [7]),
        .Q(\sr_reg[14] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [8]),
        .Q(\sr_reg[14] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[14][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[13] [9]),
        .Q(\sr_reg[14] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [0]),
        .Q(\sr_reg[1] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\sr_reg[0] [10]),
        .Q(\sr_reg[1] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [11]),
        .Q(\sr_reg[1] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [1]),
        .Q(\sr_reg[1] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [2]),
        .Q(\sr_reg[1] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [3]),
        .Q(\sr_reg[1] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [4]),
        .Q(\sr_reg[1] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [5]),
        .Q(\sr_reg[1] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [6]),
        .Q(\sr_reg[1] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [7]),
        .Q(\sr_reg[1] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [8]),
        .Q(\sr_reg[1] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[1][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\sr_reg[0] [9]),
        .Q(\sr_reg[1] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [0]),
        .Q(\sr_reg[2] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [10]),
        .Q(\sr_reg[2] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [11]),
        .Q(\sr_reg[2] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [1]),
        .Q(\sr_reg[2] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [2]),
        .Q(\sr_reg[2] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [3]),
        .Q(\sr_reg[2] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[1] [4]),
        .Q(\sr_reg[2] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[1] [5]),
        .Q(\sr_reg[2] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[1] [6]),
        .Q(\sr_reg[2] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[1] [7]),
        .Q(\sr_reg[2] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [8]),
        .Q(\sr_reg[2] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[2][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[1] [9]),
        .Q(\sr_reg[2] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [0]),
        .Q(\sr_reg[3] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [10]),
        .Q(\sr_reg[3] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [11]),
        .Q(\sr_reg[3] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [1]),
        .Q(\sr_reg[3] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [2]),
        .Q(\sr_reg[3] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [3]),
        .Q(\sr_reg[3] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[2] [4]),
        .Q(\sr_reg[3] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[2] [5]),
        .Q(\sr_reg[3] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[2] [6]),
        .Q(\sr_reg[3] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[2] [7]),
        .Q(\sr_reg[3] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [8]),
        .Q(\sr_reg[3] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[3][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[2] [9]),
        .Q(\sr_reg[3] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [0]),
        .Q(\sr_reg[4] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[3] [10]),
        .Q(\sr_reg[4] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[3] [11]),
        .Q(\sr_reg[4] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [1]),
        .Q(\sr_reg[4] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [2]),
        .Q(\sr_reg[4] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [3]),
        .Q(\sr_reg[4] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [4]),
        .Q(\sr_reg[4] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [5]),
        .Q(\sr_reg[4] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [6]),
        .Q(\sr_reg[4] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[3] [7]),
        .Q(\sr_reg[4] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[3] [8]),
        .Q(\sr_reg[4] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[4][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[3] [9]),
        .Q(\sr_reg[4] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [0]),
        .Q(\sr_reg[5] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[4] [10]),
        .Q(\sr_reg[5] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[4] [11]),
        .Q(\sr_reg[5] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [1]),
        .Q(\sr_reg[5] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [2]),
        .Q(\sr_reg[5] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [3]),
        .Q(\sr_reg[5] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [4]),
        .Q(\sr_reg[5] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [5]),
        .Q(\sr_reg[5] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [6]),
        .Q(\sr_reg[5] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[4] [7]),
        .Q(\sr_reg[5] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[4] [8]),
        .Q(\sr_reg[5] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[5][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[4] [9]),
        .Q(\sr_reg[5] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [0]),
        .Q(\sr_reg[6] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[5] [10]),
        .Q(\sr_reg[6] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[5] [11]),
        .Q(\sr_reg[6] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [1]),
        .Q(\sr_reg[6] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [2]),
        .Q(\sr_reg[6] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [3]),
        .Q(\sr_reg[6] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [4]),
        .Q(\sr_reg[6] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [5]),
        .Q(\sr_reg[6] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [6]),
        .Q(\sr_reg[6] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[5] [7]),
        .Q(\sr_reg[6] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[5] [8]),
        .Q(\sr_reg[6] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[6][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[5] [9]),
        .Q(\sr_reg[6] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [0]),
        .Q(\sr_reg[7] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[6] [10]),
        .Q(\sr_reg[7] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[6] [11]),
        .Q(\sr_reg[7] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [1]),
        .Q(\sr_reg[7] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [2]),
        .Q(\sr_reg[7] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [3]),
        .Q(\sr_reg[7] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [4]),
        .Q(\sr_reg[7] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [5]),
        .Q(\sr_reg[7] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [6]),
        .Q(\sr_reg[7] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[6] [7]),
        .Q(\sr_reg[7] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[6] [8]),
        .Q(\sr_reg[7] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[7][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[6] [9]),
        .Q(\sr_reg[7] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [0]),
        .Q(\sr_reg[8] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[7] [10]),
        .Q(\sr_reg[8] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[7] [11]),
        .Q(\sr_reg[8] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [1]),
        .Q(\sr_reg[8] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [2]),
        .Q(\sr_reg[8] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [3]),
        .Q(\sr_reg[8] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [4]),
        .Q(\sr_reg[8] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [5]),
        .Q(\sr_reg[8] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [6]),
        .Q(\sr_reg[8] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[7] [7]),
        .Q(\sr_reg[8] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[7] [8]),
        .Q(\sr_reg[8] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[8][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[7] [9]),
        .Q(\sr_reg[8] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [0]),
        .Q(\sr_reg[9] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[8] [10]),
        .Q(\sr_reg[9] [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[8] [11]),
        .Q(\sr_reg[9] [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [1]),
        .Q(\sr_reg[9] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [2]),
        .Q(\sr_reg[9] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [3]),
        .Q(\sr_reg[9] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [4]),
        .Q(\sr_reg[9] [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [5]),
        .Q(\sr_reg[9] [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [6]),
        .Q(\sr_reg[9] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\sr_reg[8] [7]),
        .Q(\sr_reg[9] [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[8] [8]),
        .Q(\sr_reg[9] [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_4/sr_reg[9][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\sr_reg[8] [9]),
        .Q(\sr_reg[9] [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/multOp 
       (.A({\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_5 ,\I_5/multOp_i_1_n_6 ,\I_5/multOp_i_1_n_7 ,\I_5/multOp_i_2_n_4 ,\I_5/multOp_i_2_n_5 ,\I_5/multOp_i_2_n_6 ,\I_5/multOp_i_2_n_7 ,\I_5/multOp_i_3_n_4 ,\I_5/multOp_i_3_n_5 ,\I_5/multOp_i_3_n_6 ,\I_5/multOp_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .PCOUT({\I_5/multOp_n_106 ,\I_5/multOp_n_107 ,\I_5/multOp_n_108 ,\I_5/multOp_n_109 ,\I_5/multOp_n_110 ,\I_5/multOp_n_111 ,\I_5/multOp_n_112 ,\I_5/multOp_n_113 ,\I_5/multOp_n_114 ,\I_5/multOp_n_115 ,\I_5/multOp_n_116 ,\I_5/multOp_n_117 ,\I_5/multOp_n_118 ,\I_5/multOp_n_119 ,\I_5/multOp_n_120 ,\I_5/multOp_n_121 ,\I_5/multOp_n_122 ,\I_5/multOp_n_123 ,\I_5/multOp_n_124 ,\I_5/multOp_n_125 ,\I_5/multOp_n_126 ,\I_5/multOp_n_127 ,\I_5/multOp_n_128 ,\I_5/multOp_n_129 ,\I_5/multOp_n_130 ,\I_5/multOp_n_131 ,\I_5/multOp_n_132 ,\I_5/multOp_n_133 ,\I_5/multOp_n_134 ,\I_5/multOp_n_135 ,\I_5/multOp_n_136 ,\I_5/multOp_n_137 ,\I_5/multOp_n_138 ,\I_5/multOp_n_139 ,\I_5/multOp_n_140 ,\I_5/multOp_n_141 ,\I_5/multOp_n_142 ,\I_5/multOp_n_143 ,\I_5/multOp_n_144 ,\I_5/multOp_n_145 ,\I_5/multOp_n_146 ,\I_5/multOp_n_147 ,\I_5/multOp_n_148 ,\I_5/multOp_n_149 ,\I_5/multOp_n_150 ,\I_5/multOp_n_151 ,\I_5/multOp_n_152 ,\I_5/multOp_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp__39_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/multOp__39_carry_n_0 ,\I_5/multOp__39_carry_n_1 ,\I_5/multOp__39_carry_n_2 ,\I_5/multOp__39_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry_i_1_n_0,multOp__39_carry_i_2_n_0,multOp__39_carry_i_3_n_0,\<const0>__0__0 }),
        .O({\I_5/multOp__39_carry_n_4 ,\I_5/multOp__39_carry_n_5 ,\I_5/multOp__39_carry_n_6 ,\I_5/multOp__39_carry_n_7 }),
        .S({multOp__39_carry_i_4_n_0,multOp__39_carry_i_5_n_0,multOp__39_carry_i_6_n_0,multOp__39_carry_i_7_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp__39_carry__0 
       (.CI(\I_5/multOp__39_carry_n_0 ),
        .CO({\I_5/multOp__39_carry__0_n_0 ,\I_5/multOp__39_carry__0_n_1 ,\I_5/multOp__39_carry__0_n_2 ,\I_5/multOp__39_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry__0_i_1_n_0,multOp__39_carry__0_i_2_n_0,multOp__39_carry__0_i_3_n_0,multOp__39_carry__0_i_4_n_0}),
        .O({\I_5/multOp__39_carry__0_n_4 ,\I_5/multOp__39_carry__0_n_5 ,\I_5/multOp__39_carry__0_n_6 ,\I_5/multOp__39_carry__0_n_7 }),
        .S({multOp__39_carry__0_i_5_n_0,multOp__39_carry__0_i_6_n_0,multOp__39_carry__0_i_7_n_0,multOp__39_carry__0_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp__39_carry__1 
       (.CI(\I_5/multOp__39_carry__0_n_0 ),
        .CO({\I_5/multOp__39_carry__1_n_0 ,\I_5/multOp__39_carry__1_n_1 ,\I_5/multOp__39_carry__1_n_2 ,\I_5/multOp__39_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({multOp__39_carry__1_i_1_n_0,multOp__39_carry__1_i_2_n_0,multOp__39_carry__1_i_3_n_0,multOp__39_carry__1_i_4_n_0}),
        .O({\I_5/multOp__39_carry__1_n_4 ,\I_5/multOp__39_carry__1_n_5 ,\I_5/multOp__39_carry__1_n_6 ,\I_5/multOp__39_carry__1_n_7 }),
        .S({multOp__39_carry__1_i_5_n_0,multOp__39_carry__1_i_6_n_0,multOp__39_carry__1_i_7_n_0,multOp__39_carry__1_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp__39_carry__2 
       (.CI(\I_5/multOp__39_carry__1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\I_5/multOp__39_carry__2_n_4 ,\I_5/multOp__39_carry__2_n_5 ,\I_5/multOp__39_carry__2_n_6 ,\I_5/multOp__39_carry__2_n_7 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,multOp__39_carry__2_i_1_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/multOp_carry_n_0 ,\I_5/multOp_carry_n_1 ,\I_5/multOp_carry_n_2 ,\I_5/multOp_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/plusOp_inferred__6_carry_n_6 ,\I_5/plusOp_inferred__6_carry_n_7 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\I_5/multOp_carry_n_4 ,\I_5/multOp_carry_n_5 ,\I_5/multOp_carry_n_6 ,\I_5/multOp_carry_n_7 }),
        .S({multOp_carry_i_1_n_0,multOp_carry_i_2_n_0,multOp_carry_i_3_n_0,\I_5/plusOp_inferred__6_carry_n_7 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_carry__0 
       (.CI(\I_5/multOp_carry_n_0 ),
        .CO({\I_5/multOp_carry__0_n_0 ,\I_5/multOp_carry__0_n_1 ,\I_5/multOp_carry__0_n_2 ,\I_5/multOp_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/plusOp_inferred__6_carry__0_n_6 ,\I_5/plusOp_inferred__6_carry__0_n_7 ,\I_5/plusOp_inferred__6_carry_n_4 ,\I_5/plusOp_inferred__6_carry_n_5 }),
        .O({\I_5/multOp_carry__0_n_4 ,\I_5/multOp_carry__0_n_5 ,\I_5/multOp_carry__0_n_6 ,\I_5/multOp_carry__0_n_7 }),
        .S({multOp_carry__0_i_1_n_0,multOp_carry__0_i_2_n_0,multOp_carry__0_i_3_n_0,multOp_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_carry__1 
       (.CI(\I_5/multOp_carry__0_n_0 ),
        .CO({\I_5/multOp_carry__1_n_0 ,\I_5/multOp_carry__1_n_1 ,\I_5/multOp_carry__1_n_2 ,\I_5/multOp_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/plusOp_inferred__6_carry__1_n_6 ,\I_5/plusOp_inferred__6_carry__1_n_7 ,\I_5/plusOp_inferred__6_carry__0_n_4 ,\I_5/plusOp_inferred__6_carry__0_n_5 }),
        .O({\I_5/multOp_carry__1_n_4 ,\I_5/multOp_carry__1_n_5 ,\I_5/multOp_carry__1_n_6 ,\I_5/multOp_carry__1_n_7 }),
        .S({multOp_carry__1_i_1_n_0,multOp_carry__1_i_2_n_0,multOp_carry__1_i_3_n_0,multOp_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_carry__2 
       (.CI(\I_5/multOp_carry__1_n_0 ),
        .CO({\I_5/multOp_carry__2_n_0 ,\I_5/multOp_carry__2_n_1 ,\I_5/multOp_carry__2_n_2 ,\I_5/multOp_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_5/plusOp_inferred__6_carry__1_n_5 }),
        .O({\I_5/multOp_carry__2_n_4 ,\I_5/multOp_carry__2_n_5 ,\I_5/multOp_carry__2_n_6 ,\I_5/multOp_carry__2_n_7 }),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,multOp_carry__2_i_1_n_0,multOp_carry__2_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_i_1 
       (.CI(\I_5/multOp_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[6][10] ,\I_5/sr_reg_n_0_[6][9] ,\I_5/sr_reg_n_0_[6][8] }),
        .O({\I_5/multOp_i_1_n_4 ,\I_5/multOp_i_1_n_5 ,\I_5/multOp_i_1_n_6 ,\I_5/multOp_i_1_n_7 }),
        .S({\I_5/multOp_i_4_n_0 ,\I_5/multOp_i_5_n_0 ,\I_5/multOp_i_6_n_0 ,\I_5/multOp_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_10 
       (.I0(\I_5/sr_reg_n_0_[6][5] ),
        .I1(\I_5/sr_reg_n_0_[7][5] ),
        .O(\I_5/multOp_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_11 
       (.I0(\I_5/sr_reg_n_0_[6][4] ),
        .I1(\I_5/sr_reg_n_0_[7][4] ),
        .O(\I_5/multOp_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_12 
       (.I0(\I_5/sr_reg_n_0_[6][3] ),
        .I1(\I_5/sr_reg_n_0_[7][3] ),
        .O(\I_5/multOp_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_13 
       (.I0(\I_5/sr_reg_n_0_[6][2] ),
        .I1(\I_5/sr_reg_n_0_[7][2] ),
        .O(\I_5/multOp_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_14 
       (.I0(\I_5/sr_reg_n_0_[6][1] ),
        .I1(\I_5/sr_reg_n_0_[7][1] ),
        .O(\I_5/multOp_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_15 
       (.I0(\I_5/sr_reg_n_0_[6][0] ),
        .I1(\I_5/sr_reg_n_0_[7][0] ),
        .O(\I_5/multOp_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_i_2 
       (.CI(\I_5/multOp_i_3_n_0 ),
        .CO({\I_5/multOp_i_2_n_0 ,\I_5/multOp_i_2_n_1 ,\I_5/multOp_i_2_n_2 ,\I_5/multOp_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[6][7] ,\I_5/sr_reg_n_0_[6][6] ,\I_5/sr_reg_n_0_[6][5] ,\I_5/sr_reg_n_0_[6][4] }),
        .O({\I_5/multOp_i_2_n_4 ,\I_5/multOp_i_2_n_5 ,\I_5/multOp_i_2_n_6 ,\I_5/multOp_i_2_n_7 }),
        .S({\I_5/multOp_i_8_n_0 ,\I_5/multOp_i_9_n_0 ,\I_5/multOp_i_10_n_0 ,\I_5/multOp_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/multOp_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/multOp_i_3_n_0 ,\I_5/multOp_i_3_n_1 ,\I_5/multOp_i_3_n_2 ,\I_5/multOp_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[6][3] ,\I_5/sr_reg_n_0_[6][2] ,\I_5/sr_reg_n_0_[6][1] ,\I_5/sr_reg_n_0_[6][0] }),
        .O({\I_5/multOp_i_3_n_4 ,\I_5/multOp_i_3_n_5 ,\I_5/multOp_i_3_n_6 ,\I_5/multOp_i_3_n_7 }),
        .S({\I_5/multOp_i_12_n_0 ,\I_5/multOp_i_13_n_0 ,\I_5/multOp_i_14_n_0 ,\I_5/multOp_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_4 
       (.I0(\I_5/sr_reg_n_0_[6][11] ),
        .I1(\I_5/sr_reg_n_0_[7][11] ),
        .O(\I_5/multOp_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_5 
       (.I0(\I_5/sr_reg_n_0_[6][10] ),
        .I1(\I_5/sr_reg_n_0_[7][10] ),
        .O(\I_5/multOp_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_6 
       (.I0(\I_5/sr_reg_n_0_[6][9] ),
        .I1(\I_5/sr_reg_n_0_[7][9] ),
        .O(\I_5/multOp_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_7 
       (.I0(\I_5/sr_reg_n_0_[6][8] ),
        .I1(\I_5/sr_reg_n_0_[7][8] ),
        .O(\I_5/multOp_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_8 
       (.I0(\I_5/sr_reg_n_0_[6][7] ),
        .I1(\I_5/sr_reg_n_0_[7][7] ),
        .O(\I_5/multOp_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/multOp_i_9 
       (.I0(\I_5/sr_reg_n_0_[6][6] ),
        .I1(\I_5/sr_reg_n_0_[7][6] ),
        .O(\I_5/multOp_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__1_n_4 ),
        .Q(\I_5/output_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__4_n_6 ),
        .Q(\I_5/output_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__4_n_5 ),
        .Q(\I_5/output_reg_n_0_[11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__2_n_7 ),
        .Q(\I_5/output_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__2_n_6 ),
        .Q(\I_5/output_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__2_n_5 ),
        .Q(\I_5/output_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__2_n_4 ),
        .Q(\I_5/output_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__3_n_7 ),
        .Q(\I_5/output_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__3_n_6 ),
        .Q(\I_5/output_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__3_n_5 ),
        .Q(\I_5/output_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__3_n_4 ),
        .Q(\I_5/output_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/output_reg[9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_phase_i_2_n_0),
        .D(\I_5/plusOp_inferred__7__62_carry__4_n_7 ),
        .Q(\I_5/output_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/plusOp 
       (.A({\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_5 ,\I_5/plusOp_inferred__3_carry__1_n_6 ,\I_5/plusOp_inferred__3_carry__1_n_7 ,\I_5/plusOp_inferred__3_carry__0_n_4 ,\I_5/plusOp_inferred__3_carry__0_n_5 ,\I_5/plusOp_inferred__3_carry__0_n_6 ,\I_5/plusOp_inferred__3_carry__0_n_7 ,\I_5/plusOp_inferred__3_carry_n_4 ,\I_5/plusOp_inferred__3_carry_n_5 ,\I_5/plusOp_inferred__3_carry_n_6 ,\I_5/plusOp_inferred__3_carry_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_5/multOp_n_106 ,\I_5/multOp_n_107 ,\I_5/multOp_n_108 ,\I_5/multOp_n_109 ,\I_5/multOp_n_110 ,\I_5/multOp_n_111 ,\I_5/multOp_n_112 ,\I_5/multOp_n_113 ,\I_5/multOp_n_114 ,\I_5/multOp_n_115 ,\I_5/multOp_n_116 ,\I_5/multOp_n_117 ,\I_5/multOp_n_118 ,\I_5/multOp_n_119 ,\I_5/multOp_n_120 ,\I_5/multOp_n_121 ,\I_5/multOp_n_122 ,\I_5/multOp_n_123 ,\I_5/multOp_n_124 ,\I_5/multOp_n_125 ,\I_5/multOp_n_126 ,\I_5/multOp_n_127 ,\I_5/multOp_n_128 ,\I_5/multOp_n_129 ,\I_5/multOp_n_130 ,\I_5/multOp_n_131 ,\I_5/multOp_n_132 ,\I_5/multOp_n_133 ,\I_5/multOp_n_134 ,\I_5/multOp_n_135 ,\I_5/multOp_n_136 ,\I_5/multOp_n_137 ,\I_5/multOp_n_138 ,\I_5/multOp_n_139 ,\I_5/multOp_n_140 ,\I_5/multOp_n_141 ,\I_5/multOp_n_142 ,\I_5/multOp_n_143 ,\I_5/multOp_n_144 ,\I_5/multOp_n_145 ,\I_5/multOp_n_146 ,\I_5/multOp_n_147 ,\I_5/multOp_n_148 ,\I_5/multOp_n_149 ,\I_5/multOp_n_150 ,\I_5/multOp_n_151 ,\I_5/multOp_n_152 ,\I_5/multOp_n_153 }),
        .PCOUT({\I_5/plusOp_n_106 ,\I_5/plusOp_n_107 ,\I_5/plusOp_n_108 ,\I_5/plusOp_n_109 ,\I_5/plusOp_n_110 ,\I_5/plusOp_n_111 ,\I_5/plusOp_n_112 ,\I_5/plusOp_n_113 ,\I_5/plusOp_n_114 ,\I_5/plusOp_n_115 ,\I_5/plusOp_n_116 ,\I_5/plusOp_n_117 ,\I_5/plusOp_n_118 ,\I_5/plusOp_n_119 ,\I_5/plusOp_n_120 ,\I_5/plusOp_n_121 ,\I_5/plusOp_n_122 ,\I_5/plusOp_n_123 ,\I_5/plusOp_n_124 ,\I_5/plusOp_n_125 ,\I_5/plusOp_n_126 ,\I_5/plusOp_n_127 ,\I_5/plusOp_n_128 ,\I_5/plusOp_n_129 ,\I_5/plusOp_n_130 ,\I_5/plusOp_n_131 ,\I_5/plusOp_n_132 ,\I_5/plusOp_n_133 ,\I_5/plusOp_n_134 ,\I_5/plusOp_n_135 ,\I_5/plusOp_n_136 ,\I_5/plusOp_n_137 ,\I_5/plusOp_n_138 ,\I_5/plusOp_n_139 ,\I_5/plusOp_n_140 ,\I_5/plusOp_n_141 ,\I_5/plusOp_n_142 ,\I_5/plusOp_n_143 ,\I_5/plusOp_n_144 ,\I_5/plusOp_n_145 ,\I_5/plusOp_n_146 ,\I_5/plusOp_n_147 ,\I_5/plusOp_n_148 ,\I_5/plusOp_n_149 ,\I_5/plusOp_n_150 ,\I_5/plusOp_n_151 ,\I_5/plusOp_n_152 ,\I_5/plusOp_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/plusOp__0 
       (.A({\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_5 ,\I_5/plusOp__0_i_1_n_6 ,\I_5/plusOp__0_i_1_n_7 ,\I_5/plusOp__0_i_2_n_4 ,\I_5/plusOp__0_i_2_n_5 ,\I_5/plusOp__0_i_2_n_6 ,\I_5/plusOp__0_i_2_n_7 ,\I_5/plusOp__0_i_3_n_4 ,\I_5/plusOp__0_i_3_n_5 ,\I_5/plusOp__0_i_3_n_6 ,\I_5/plusOp__0_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_5/plusOp_n_106 ,\I_5/plusOp_n_107 ,\I_5/plusOp_n_108 ,\I_5/plusOp_n_109 ,\I_5/plusOp_n_110 ,\I_5/plusOp_n_111 ,\I_5/plusOp_n_112 ,\I_5/plusOp_n_113 ,\I_5/plusOp_n_114 ,\I_5/plusOp_n_115 ,\I_5/plusOp_n_116 ,\I_5/plusOp_n_117 ,\I_5/plusOp_n_118 ,\I_5/plusOp_n_119 ,\I_5/plusOp_n_120 ,\I_5/plusOp_n_121 ,\I_5/plusOp_n_122 ,\I_5/plusOp_n_123 ,\I_5/plusOp_n_124 ,\I_5/plusOp_n_125 ,\I_5/plusOp_n_126 ,\I_5/plusOp_n_127 ,\I_5/plusOp_n_128 ,\I_5/plusOp_n_129 ,\I_5/plusOp_n_130 ,\I_5/plusOp_n_131 ,\I_5/plusOp_n_132 ,\I_5/plusOp_n_133 ,\I_5/plusOp_n_134 ,\I_5/plusOp_n_135 ,\I_5/plusOp_n_136 ,\I_5/plusOp_n_137 ,\I_5/plusOp_n_138 ,\I_5/plusOp_n_139 ,\I_5/plusOp_n_140 ,\I_5/plusOp_n_141 ,\I_5/plusOp_n_142 ,\I_5/plusOp_n_143 ,\I_5/plusOp_n_144 ,\I_5/plusOp_n_145 ,\I_5/plusOp_n_146 ,\I_5/plusOp_n_147 ,\I_5/plusOp_n_148 ,\I_5/plusOp_n_149 ,\I_5/plusOp_n_150 ,\I_5/plusOp_n_151 ,\I_5/plusOp_n_152 ,\I_5/plusOp_n_153 }),
        .PCOUT({\I_5/plusOp__0_n_106 ,\I_5/plusOp__0_n_107 ,\I_5/plusOp__0_n_108 ,\I_5/plusOp__0_n_109 ,\I_5/plusOp__0_n_110 ,\I_5/plusOp__0_n_111 ,\I_5/plusOp__0_n_112 ,\I_5/plusOp__0_n_113 ,\I_5/plusOp__0_n_114 ,\I_5/plusOp__0_n_115 ,\I_5/plusOp__0_n_116 ,\I_5/plusOp__0_n_117 ,\I_5/plusOp__0_n_118 ,\I_5/plusOp__0_n_119 ,\I_5/plusOp__0_n_120 ,\I_5/plusOp__0_n_121 ,\I_5/plusOp__0_n_122 ,\I_5/plusOp__0_n_123 ,\I_5/plusOp__0_n_124 ,\I_5/plusOp__0_n_125 ,\I_5/plusOp__0_n_126 ,\I_5/plusOp__0_n_127 ,\I_5/plusOp__0_n_128 ,\I_5/plusOp__0_n_129 ,\I_5/plusOp__0_n_130 ,\I_5/plusOp__0_n_131 ,\I_5/plusOp__0_n_132 ,\I_5/plusOp__0_n_133 ,\I_5/plusOp__0_n_134 ,\I_5/plusOp__0_n_135 ,\I_5/plusOp__0_n_136 ,\I_5/plusOp__0_n_137 ,\I_5/plusOp__0_n_138 ,\I_5/plusOp__0_n_139 ,\I_5/plusOp__0_n_140 ,\I_5/plusOp__0_n_141 ,\I_5/plusOp__0_n_142 ,\I_5/plusOp__0_n_143 ,\I_5/plusOp__0_n_144 ,\I_5/plusOp__0_n_145 ,\I_5/plusOp__0_n_146 ,\I_5/plusOp__0_n_147 ,\I_5/plusOp__0_n_148 ,\I_5/plusOp__0_n_149 ,\I_5/plusOp__0_n_150 ,\I_5/plusOp__0_n_151 ,\I_5/plusOp__0_n_152 ,\I_5/plusOp__0_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__0_i_1 
       (.CI(\I_5/plusOp__0_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[5][10] ,\I_5/sr_reg_n_0_[5][9] ,\I_5/sr_reg_n_0_[5][8] }),
        .O({\I_5/plusOp__0_i_1_n_4 ,\I_5/plusOp__0_i_1_n_5 ,\I_5/plusOp__0_i_1_n_6 ,\I_5/plusOp__0_i_1_n_7 }),
        .S({\I_5/plusOp__0_i_4_n_0 ,\I_5/plusOp__0_i_5_n_0 ,\I_5/plusOp__0_i_6_n_0 ,\I_5/plusOp__0_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_10 
       (.I0(\I_5/sr_reg_n_0_[5][5] ),
        .I1(\I_5/sr_reg_n_0_[8][5] ),
        .O(\I_5/plusOp__0_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_11 
       (.I0(\I_5/sr_reg_n_0_[5][4] ),
        .I1(\I_5/sr_reg_n_0_[8][4] ),
        .O(\I_5/plusOp__0_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_12 
       (.I0(\I_5/sr_reg_n_0_[5][3] ),
        .I1(\I_5/sr_reg_n_0_[8][3] ),
        .O(\I_5/plusOp__0_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_13 
       (.I0(\I_5/sr_reg_n_0_[5][2] ),
        .I1(\I_5/sr_reg_n_0_[8][2] ),
        .O(\I_5/plusOp__0_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_14 
       (.I0(\I_5/sr_reg_n_0_[5][1] ),
        .I1(\I_5/sr_reg_n_0_[8][1] ),
        .O(\I_5/plusOp__0_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_15 
       (.I0(\I_5/sr_reg_n_0_[5][0] ),
        .I1(\I_5/sr_reg_n_0_[8][0] ),
        .O(\I_5/plusOp__0_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__0_i_2 
       (.CI(\I_5/plusOp__0_i_3_n_0 ),
        .CO({\I_5/plusOp__0_i_2_n_0 ,\I_5/plusOp__0_i_2_n_1 ,\I_5/plusOp__0_i_2_n_2 ,\I_5/plusOp__0_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[5][7] ,\I_5/sr_reg_n_0_[5][6] ,\I_5/sr_reg_n_0_[5][5] ,\I_5/sr_reg_n_0_[5][4] }),
        .O({\I_5/plusOp__0_i_2_n_4 ,\I_5/plusOp__0_i_2_n_5 ,\I_5/plusOp__0_i_2_n_6 ,\I_5/plusOp__0_i_2_n_7 }),
        .S({\I_5/plusOp__0_i_8_n_0 ,\I_5/plusOp__0_i_9_n_0 ,\I_5/plusOp__0_i_10_n_0 ,\I_5/plusOp__0_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__0_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp__0_i_3_n_0 ,\I_5/plusOp__0_i_3_n_1 ,\I_5/plusOp__0_i_3_n_2 ,\I_5/plusOp__0_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[5][3] ,\I_5/sr_reg_n_0_[5][2] ,\I_5/sr_reg_n_0_[5][1] ,\I_5/sr_reg_n_0_[5][0] }),
        .O({\I_5/plusOp__0_i_3_n_4 ,\I_5/plusOp__0_i_3_n_5 ,\I_5/plusOp__0_i_3_n_6 ,\I_5/plusOp__0_i_3_n_7 }),
        .S({\I_5/plusOp__0_i_12_n_0 ,\I_5/plusOp__0_i_13_n_0 ,\I_5/plusOp__0_i_14_n_0 ,\I_5/plusOp__0_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_4 
       (.I0(\I_5/sr_reg_n_0_[5][11] ),
        .I1(\I_5/sr_reg_n_0_[8][11] ),
        .O(\I_5/plusOp__0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_5 
       (.I0(\I_5/sr_reg_n_0_[5][10] ),
        .I1(\I_5/sr_reg_n_0_[8][10] ),
        .O(\I_5/plusOp__0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_6 
       (.I0(\I_5/sr_reg_n_0_[5][9] ),
        .I1(\I_5/sr_reg_n_0_[8][9] ),
        .O(\I_5/plusOp__0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_7 
       (.I0(\I_5/sr_reg_n_0_[5][8] ),
        .I1(\I_5/sr_reg_n_0_[8][8] ),
        .O(\I_5/plusOp__0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_8 
       (.I0(\I_5/sr_reg_n_0_[5][7] ),
        .I1(\I_5/sr_reg_n_0_[8][7] ),
        .O(\I_5/plusOp__0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__0_i_9 
       (.I0(\I_5/sr_reg_n_0_[5][6] ),
        .I1(\I_5/sr_reg_n_0_[8][6] ),
        .O(\I_5/plusOp__0_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/plusOp__1 
       (.A({\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_5 ,\I_5/plusOp__1_i_1_n_6 ,\I_5/plusOp__1_i_1_n_7 ,\I_5/plusOp__1_i_2_n_4 ,\I_5/plusOp__1_i_2_n_5 ,\I_5/plusOp__1_i_2_n_6 ,\I_5/plusOp__1_i_2_n_7 ,\I_5/plusOp__1_i_3_n_4 ,\I_5/plusOp__1_i_3_n_5 ,\I_5/plusOp__1_i_3_n_6 ,\I_5/plusOp__1_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_5/plusOp__0_n_106 ,\I_5/plusOp__0_n_107 ,\I_5/plusOp__0_n_108 ,\I_5/plusOp__0_n_109 ,\I_5/plusOp__0_n_110 ,\I_5/plusOp__0_n_111 ,\I_5/plusOp__0_n_112 ,\I_5/plusOp__0_n_113 ,\I_5/plusOp__0_n_114 ,\I_5/plusOp__0_n_115 ,\I_5/plusOp__0_n_116 ,\I_5/plusOp__0_n_117 ,\I_5/plusOp__0_n_118 ,\I_5/plusOp__0_n_119 ,\I_5/plusOp__0_n_120 ,\I_5/plusOp__0_n_121 ,\I_5/plusOp__0_n_122 ,\I_5/plusOp__0_n_123 ,\I_5/plusOp__0_n_124 ,\I_5/plusOp__0_n_125 ,\I_5/plusOp__0_n_126 ,\I_5/plusOp__0_n_127 ,\I_5/plusOp__0_n_128 ,\I_5/plusOp__0_n_129 ,\I_5/plusOp__0_n_130 ,\I_5/plusOp__0_n_131 ,\I_5/plusOp__0_n_132 ,\I_5/plusOp__0_n_133 ,\I_5/plusOp__0_n_134 ,\I_5/plusOp__0_n_135 ,\I_5/plusOp__0_n_136 ,\I_5/plusOp__0_n_137 ,\I_5/plusOp__0_n_138 ,\I_5/plusOp__0_n_139 ,\I_5/plusOp__0_n_140 ,\I_5/plusOp__0_n_141 ,\I_5/plusOp__0_n_142 ,\I_5/plusOp__0_n_143 ,\I_5/plusOp__0_n_144 ,\I_5/plusOp__0_n_145 ,\I_5/plusOp__0_n_146 ,\I_5/plusOp__0_n_147 ,\I_5/plusOp__0_n_148 ,\I_5/plusOp__0_n_149 ,\I_5/plusOp__0_n_150 ,\I_5/plusOp__0_n_151 ,\I_5/plusOp__0_n_152 ,\I_5/plusOp__0_n_153 }),
        .PCOUT({\I_5/plusOp__1_n_106 ,\I_5/plusOp__1_n_107 ,\I_5/plusOp__1_n_108 ,\I_5/plusOp__1_n_109 ,\I_5/plusOp__1_n_110 ,\I_5/plusOp__1_n_111 ,\I_5/plusOp__1_n_112 ,\I_5/plusOp__1_n_113 ,\I_5/plusOp__1_n_114 ,\I_5/plusOp__1_n_115 ,\I_5/plusOp__1_n_116 ,\I_5/plusOp__1_n_117 ,\I_5/plusOp__1_n_118 ,\I_5/plusOp__1_n_119 ,\I_5/plusOp__1_n_120 ,\I_5/plusOp__1_n_121 ,\I_5/plusOp__1_n_122 ,\I_5/plusOp__1_n_123 ,\I_5/plusOp__1_n_124 ,\I_5/plusOp__1_n_125 ,\I_5/plusOp__1_n_126 ,\I_5/plusOp__1_n_127 ,\I_5/plusOp__1_n_128 ,\I_5/plusOp__1_n_129 ,\I_5/plusOp__1_n_130 ,\I_5/plusOp__1_n_131 ,\I_5/plusOp__1_n_132 ,\I_5/plusOp__1_n_133 ,\I_5/plusOp__1_n_134 ,\I_5/plusOp__1_n_135 ,\I_5/plusOp__1_n_136 ,\I_5/plusOp__1_n_137 ,\I_5/plusOp__1_n_138 ,\I_5/plusOp__1_n_139 ,\I_5/plusOp__1_n_140 ,\I_5/plusOp__1_n_141 ,\I_5/plusOp__1_n_142 ,\I_5/plusOp__1_n_143 ,\I_5/plusOp__1_n_144 ,\I_5/plusOp__1_n_145 ,\I_5/plusOp__1_n_146 ,\I_5/plusOp__1_n_147 ,\I_5/plusOp__1_n_148 ,\I_5/plusOp__1_n_149 ,\I_5/plusOp__1_n_150 ,\I_5/plusOp__1_n_151 ,\I_5/plusOp__1_n_152 ,\I_5/plusOp__1_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__1_i_1 
       (.CI(\I_5/plusOp__1_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[4][10] ,\I_5/sr_reg_n_0_[4][9] ,\I_5/sr_reg_n_0_[4][8] }),
        .O({\I_5/plusOp__1_i_1_n_4 ,\I_5/plusOp__1_i_1_n_5 ,\I_5/plusOp__1_i_1_n_6 ,\I_5/plusOp__1_i_1_n_7 }),
        .S({\I_5/plusOp__1_i_4_n_0 ,\I_5/plusOp__1_i_5_n_0 ,\I_5/plusOp__1_i_6_n_0 ,\I_5/plusOp__1_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_10 
       (.I0(\I_5/sr_reg_n_0_[4][5] ),
        .I1(\I_5/sr_reg_n_0_[9][5] ),
        .O(\I_5/plusOp__1_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_11 
       (.I0(\I_5/sr_reg_n_0_[4][4] ),
        .I1(\I_5/sr_reg_n_0_[9][4] ),
        .O(\I_5/plusOp__1_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_12 
       (.I0(\I_5/sr_reg_n_0_[4][3] ),
        .I1(\I_5/sr_reg_n_0_[9][3] ),
        .O(\I_5/plusOp__1_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_13 
       (.I0(\I_5/sr_reg_n_0_[4][2] ),
        .I1(\I_5/sr_reg_n_0_[9][2] ),
        .O(\I_5/plusOp__1_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_14 
       (.I0(\I_5/sr_reg_n_0_[4][1] ),
        .I1(\I_5/sr_reg_n_0_[9][1] ),
        .O(\I_5/plusOp__1_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_15 
       (.I0(\I_5/sr_reg_n_0_[4][0] ),
        .I1(\I_5/sr_reg_n_0_[9][0] ),
        .O(\I_5/plusOp__1_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__1_i_2 
       (.CI(\I_5/plusOp__1_i_3_n_0 ),
        .CO({\I_5/plusOp__1_i_2_n_0 ,\I_5/plusOp__1_i_2_n_1 ,\I_5/plusOp__1_i_2_n_2 ,\I_5/plusOp__1_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[4][7] ,\I_5/sr_reg_n_0_[4][6] ,\I_5/sr_reg_n_0_[4][5] ,\I_5/sr_reg_n_0_[4][4] }),
        .O({\I_5/plusOp__1_i_2_n_4 ,\I_5/plusOp__1_i_2_n_5 ,\I_5/plusOp__1_i_2_n_6 ,\I_5/plusOp__1_i_2_n_7 }),
        .S({\I_5/plusOp__1_i_8_n_0 ,\I_5/plusOp__1_i_9_n_0 ,\I_5/plusOp__1_i_10_n_0 ,\I_5/plusOp__1_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__1_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp__1_i_3_n_0 ,\I_5/plusOp__1_i_3_n_1 ,\I_5/plusOp__1_i_3_n_2 ,\I_5/plusOp__1_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[4][3] ,\I_5/sr_reg_n_0_[4][2] ,\I_5/sr_reg_n_0_[4][1] ,\I_5/sr_reg_n_0_[4][0] }),
        .O({\I_5/plusOp__1_i_3_n_4 ,\I_5/plusOp__1_i_3_n_5 ,\I_5/plusOp__1_i_3_n_6 ,\I_5/plusOp__1_i_3_n_7 }),
        .S({\I_5/plusOp__1_i_12_n_0 ,\I_5/plusOp__1_i_13_n_0 ,\I_5/plusOp__1_i_14_n_0 ,\I_5/plusOp__1_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_4 
       (.I0(\I_5/sr_reg_n_0_[4][11] ),
        .I1(\I_5/sr_reg_n_0_[9][11] ),
        .O(\I_5/plusOp__1_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_5 
       (.I0(\I_5/sr_reg_n_0_[4][10] ),
        .I1(\I_5/sr_reg_n_0_[9][10] ),
        .O(\I_5/plusOp__1_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_6 
       (.I0(\I_5/sr_reg_n_0_[4][9] ),
        .I1(\I_5/sr_reg_n_0_[9][9] ),
        .O(\I_5/plusOp__1_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_7 
       (.I0(\I_5/sr_reg_n_0_[4][8] ),
        .I1(\I_5/sr_reg_n_0_[9][8] ),
        .O(\I_5/plusOp__1_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_8 
       (.I0(\I_5/sr_reg_n_0_[4][7] ),
        .I1(\I_5/sr_reg_n_0_[9][7] ),
        .O(\I_5/plusOp__1_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__1_i_9 
       (.I0(\I_5/sr_reg_n_0_[4][6] ),
        .I1(\I_5/sr_reg_n_0_[9][6] ),
        .O(\I_5/plusOp__1_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/plusOp__2 
       (.A({\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_5 ,\I_5/plusOp__2_i_1_n_6 ,\I_5/plusOp__2_i_1_n_7 ,\I_5/plusOp__2_i_2_n_4 ,\I_5/plusOp__2_i_2_n_5 ,\I_5/plusOp__2_i_2_n_6 ,\I_5/plusOp__2_i_2_n_7 ,\I_5/plusOp__2_i_3_n_4 ,\I_5/plusOp__2_i_3_n_5 ,\I_5/plusOp__2_i_3_n_6 ,\I_5/plusOp__2_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .PCIN({\I_5/plusOp__1_n_106 ,\I_5/plusOp__1_n_107 ,\I_5/plusOp__1_n_108 ,\I_5/plusOp__1_n_109 ,\I_5/plusOp__1_n_110 ,\I_5/plusOp__1_n_111 ,\I_5/plusOp__1_n_112 ,\I_5/plusOp__1_n_113 ,\I_5/plusOp__1_n_114 ,\I_5/plusOp__1_n_115 ,\I_5/plusOp__1_n_116 ,\I_5/plusOp__1_n_117 ,\I_5/plusOp__1_n_118 ,\I_5/plusOp__1_n_119 ,\I_5/plusOp__1_n_120 ,\I_5/plusOp__1_n_121 ,\I_5/plusOp__1_n_122 ,\I_5/plusOp__1_n_123 ,\I_5/plusOp__1_n_124 ,\I_5/plusOp__1_n_125 ,\I_5/plusOp__1_n_126 ,\I_5/plusOp__1_n_127 ,\I_5/plusOp__1_n_128 ,\I_5/plusOp__1_n_129 ,\I_5/plusOp__1_n_130 ,\I_5/plusOp__1_n_131 ,\I_5/plusOp__1_n_132 ,\I_5/plusOp__1_n_133 ,\I_5/plusOp__1_n_134 ,\I_5/plusOp__1_n_135 ,\I_5/plusOp__1_n_136 ,\I_5/plusOp__1_n_137 ,\I_5/plusOp__1_n_138 ,\I_5/plusOp__1_n_139 ,\I_5/plusOp__1_n_140 ,\I_5/plusOp__1_n_141 ,\I_5/plusOp__1_n_142 ,\I_5/plusOp__1_n_143 ,\I_5/plusOp__1_n_144 ,\I_5/plusOp__1_n_145 ,\I_5/plusOp__1_n_146 ,\I_5/plusOp__1_n_147 ,\I_5/plusOp__1_n_148 ,\I_5/plusOp__1_n_149 ,\I_5/plusOp__1_n_150 ,\I_5/plusOp__1_n_151 ,\I_5/plusOp__1_n_152 ,\I_5/plusOp__1_n_153 }),
        .PCOUT({\I_5/plusOp__2_n_106 ,\I_5/plusOp__2_n_107 ,\I_5/plusOp__2_n_108 ,\I_5/plusOp__2_n_109 ,\I_5/plusOp__2_n_110 ,\I_5/plusOp__2_n_111 ,\I_5/plusOp__2_n_112 ,\I_5/plusOp__2_n_113 ,\I_5/plusOp__2_n_114 ,\I_5/plusOp__2_n_115 ,\I_5/plusOp__2_n_116 ,\I_5/plusOp__2_n_117 ,\I_5/plusOp__2_n_118 ,\I_5/plusOp__2_n_119 ,\I_5/plusOp__2_n_120 ,\I_5/plusOp__2_n_121 ,\I_5/plusOp__2_n_122 ,\I_5/plusOp__2_n_123 ,\I_5/plusOp__2_n_124 ,\I_5/plusOp__2_n_125 ,\I_5/plusOp__2_n_126 ,\I_5/plusOp__2_n_127 ,\I_5/plusOp__2_n_128 ,\I_5/plusOp__2_n_129 ,\I_5/plusOp__2_n_130 ,\I_5/plusOp__2_n_131 ,\I_5/plusOp__2_n_132 ,\I_5/plusOp__2_n_133 ,\I_5/plusOp__2_n_134 ,\I_5/plusOp__2_n_135 ,\I_5/plusOp__2_n_136 ,\I_5/plusOp__2_n_137 ,\I_5/plusOp__2_n_138 ,\I_5/plusOp__2_n_139 ,\I_5/plusOp__2_n_140 ,\I_5/plusOp__2_n_141 ,\I_5/plusOp__2_n_142 ,\I_5/plusOp__2_n_143 ,\I_5/plusOp__2_n_144 ,\I_5/plusOp__2_n_145 ,\I_5/plusOp__2_n_146 ,\I_5/plusOp__2_n_147 ,\I_5/plusOp__2_n_148 ,\I_5/plusOp__2_n_149 ,\I_5/plusOp__2_n_150 ,\I_5/plusOp__2_n_151 ,\I_5/plusOp__2_n_152 ,\I_5/plusOp__2_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__2_i_1 
       (.CI(\I_5/plusOp__2_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[3][10] ,\I_5/sr_reg_n_0_[3][9] ,\I_5/sr_reg_n_0_[3][8] }),
        .O({\I_5/plusOp__2_i_1_n_4 ,\I_5/plusOp__2_i_1_n_5 ,\I_5/plusOp__2_i_1_n_6 ,\I_5/plusOp__2_i_1_n_7 }),
        .S({\I_5/plusOp__2_i_4_n_0 ,\I_5/plusOp__2_i_5_n_0 ,\I_5/plusOp__2_i_6_n_0 ,\I_5/plusOp__2_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_10 
       (.I0(\I_5/sr_reg_n_0_[3][5] ),
        .I1(\I_5/sr_reg_n_0_[10][5] ),
        .O(\I_5/plusOp__2_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_11 
       (.I0(\I_5/sr_reg_n_0_[3][4] ),
        .I1(\I_5/sr_reg_n_0_[10][4] ),
        .O(\I_5/plusOp__2_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_12 
       (.I0(\I_5/sr_reg_n_0_[3][3] ),
        .I1(\I_5/sr_reg_n_0_[10][3] ),
        .O(\I_5/plusOp__2_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_13 
       (.I0(\I_5/sr_reg_n_0_[3][2] ),
        .I1(\I_5/sr_reg_n_0_[10][2] ),
        .O(\I_5/plusOp__2_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_14 
       (.I0(\I_5/sr_reg_n_0_[3][1] ),
        .I1(\I_5/sr_reg_n_0_[10][1] ),
        .O(\I_5/plusOp__2_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_15 
       (.I0(\I_5/sr_reg_n_0_[3][0] ),
        .I1(\I_5/sr_reg_n_0_[10][0] ),
        .O(\I_5/plusOp__2_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__2_i_2 
       (.CI(\I_5/plusOp__2_i_3_n_0 ),
        .CO({\I_5/plusOp__2_i_2_n_0 ,\I_5/plusOp__2_i_2_n_1 ,\I_5/plusOp__2_i_2_n_2 ,\I_5/plusOp__2_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[3][7] ,\I_5/sr_reg_n_0_[3][6] ,\I_5/sr_reg_n_0_[3][5] ,\I_5/sr_reg_n_0_[3][4] }),
        .O({\I_5/plusOp__2_i_2_n_4 ,\I_5/plusOp__2_i_2_n_5 ,\I_5/plusOp__2_i_2_n_6 ,\I_5/plusOp__2_i_2_n_7 }),
        .S({\I_5/plusOp__2_i_8_n_0 ,\I_5/plusOp__2_i_9_n_0 ,\I_5/plusOp__2_i_10_n_0 ,\I_5/plusOp__2_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__2_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp__2_i_3_n_0 ,\I_5/plusOp__2_i_3_n_1 ,\I_5/plusOp__2_i_3_n_2 ,\I_5/plusOp__2_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[3][3] ,\I_5/sr_reg_n_0_[3][2] ,\I_5/sr_reg_n_0_[3][1] ,\I_5/sr_reg_n_0_[3][0] }),
        .O({\I_5/plusOp__2_i_3_n_4 ,\I_5/plusOp__2_i_3_n_5 ,\I_5/plusOp__2_i_3_n_6 ,\I_5/plusOp__2_i_3_n_7 }),
        .S({\I_5/plusOp__2_i_12_n_0 ,\I_5/plusOp__2_i_13_n_0 ,\I_5/plusOp__2_i_14_n_0 ,\I_5/plusOp__2_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_4 
       (.I0(\I_5/sr_reg_n_0_[3][11] ),
        .I1(\I_5/sr_reg_n_0_[10][11] ),
        .O(\I_5/plusOp__2_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_5 
       (.I0(\I_5/sr_reg_n_0_[3][10] ),
        .I1(\I_5/sr_reg_n_0_[10][10] ),
        .O(\I_5/plusOp__2_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_6 
       (.I0(\I_5/sr_reg_n_0_[3][9] ),
        .I1(\I_5/sr_reg_n_0_[10][9] ),
        .O(\I_5/plusOp__2_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_7 
       (.I0(\I_5/sr_reg_n_0_[3][8] ),
        .I1(\I_5/sr_reg_n_0_[10][8] ),
        .O(\I_5/plusOp__2_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_8 
       (.I0(\I_5/sr_reg_n_0_[3][7] ),
        .I1(\I_5/sr_reg_n_0_[10][7] ),
        .O(\I_5/plusOp__2_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__2_i_9 
       (.I0(\I_5/sr_reg_n_0_[3][6] ),
        .I1(\I_5/sr_reg_n_0_[10][6] ),
        .O(\I_5/plusOp__2_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-11 {cell *THIS*}} {SYNTH-13 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(0),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    \I_5/plusOp__3 
       (.A({\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_5 ,\I_5/plusOp__3_i_1_n_6 ,\I_5/plusOp__3_i_1_n_7 ,\I_5/plusOp__3_i_2_n_4 ,\I_5/plusOp__3_i_2_n_5 ,\I_5/plusOp__3_i_2_n_6 ,\I_5/plusOp__3_i_2_n_7 ,\I_5/plusOp__3_i_3_n_4 ,\I_5/plusOp__3_i_3_n_5 ,\I_5/plusOp__3_i_3_n_6 ,\I_5/plusOp__3_i_3_n_7 }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(\<const0>__0__0 ),
        .CEP(\<const0>__0__0 ),
        .CLK(\<const0>__0__0 ),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({\I_5/plusOp__3_n_58 ,\I_5/plusOp__3_n_59 ,\I_5/plusOp__3_n_60 ,\I_5/plusOp__3_n_61 ,\I_5/plusOp__3_n_62 ,\I_5/plusOp__3_n_63 ,\I_5/plusOp__3_n_64 ,\I_5/plusOp__3_n_65 ,\I_5/plusOp__3_n_66 ,\I_5/plusOp__3_n_67 ,\I_5/plusOp__3_n_68 ,\I_5/plusOp__3_n_69 ,\I_5/plusOp__3_n_70 ,\I_5/plusOp__3_n_71 ,\I_5/plusOp__3_n_72 ,\I_5/plusOp__3_n_73 ,\I_5/plusOp__3_n_74 ,\I_5/plusOp__3_n_75 ,\I_5/plusOp__3_n_76 ,\I_5/plusOp__3_n_77 ,\I_5/plusOp__3_n_78 ,\I_5/plusOp__3_n_79 ,\I_5/plusOp__3_n_80 ,\I_5/plusOp__3_n_81 ,\I_5/plusOp__3_n_82 ,\I_5/plusOp__3_n_83 ,\I_5/plusOp__3_n_84 ,\I_5/plusOp__3_n_85 ,\I_5/plusOp__3_n_86 ,\I_5/plusOp__3_n_87 ,\I_5/plusOp__3_n_88 ,\I_5/plusOp__3_n_89 ,\I_5/plusOp__3_n_90 ,\I_5/plusOp__3_n_91 ,\I_5/plusOp__3_n_92 ,\I_5/plusOp__3_n_93 ,\I_5/plusOp__3_n_94 ,\I_5/plusOp__3_n_95 ,\I_5/plusOp__3_n_96 ,\I_5/plusOp__3_n_97 ,\I_5/plusOp__3_n_98 ,\I_5/plusOp__3_n_99 ,\I_5/plusOp__3_n_100 ,\I_5/plusOp__3_n_101 ,\I_5/plusOp__3_n_102 ,\I_5/plusOp__3_n_103 ,\I_5/plusOp__3_n_104 ,\I_5/plusOp__3_n_105 }),
        .PCIN({\I_5/plusOp__2_n_106 ,\I_5/plusOp__2_n_107 ,\I_5/plusOp__2_n_108 ,\I_5/plusOp__2_n_109 ,\I_5/plusOp__2_n_110 ,\I_5/plusOp__2_n_111 ,\I_5/plusOp__2_n_112 ,\I_5/plusOp__2_n_113 ,\I_5/plusOp__2_n_114 ,\I_5/plusOp__2_n_115 ,\I_5/plusOp__2_n_116 ,\I_5/plusOp__2_n_117 ,\I_5/plusOp__2_n_118 ,\I_5/plusOp__2_n_119 ,\I_5/plusOp__2_n_120 ,\I_5/plusOp__2_n_121 ,\I_5/plusOp__2_n_122 ,\I_5/plusOp__2_n_123 ,\I_5/plusOp__2_n_124 ,\I_5/plusOp__2_n_125 ,\I_5/plusOp__2_n_126 ,\I_5/plusOp__2_n_127 ,\I_5/plusOp__2_n_128 ,\I_5/plusOp__2_n_129 ,\I_5/plusOp__2_n_130 ,\I_5/plusOp__2_n_131 ,\I_5/plusOp__2_n_132 ,\I_5/plusOp__2_n_133 ,\I_5/plusOp__2_n_134 ,\I_5/plusOp__2_n_135 ,\I_5/plusOp__2_n_136 ,\I_5/plusOp__2_n_137 ,\I_5/plusOp__2_n_138 ,\I_5/plusOp__2_n_139 ,\I_5/plusOp__2_n_140 ,\I_5/plusOp__2_n_141 ,\I_5/plusOp__2_n_142 ,\I_5/plusOp__2_n_143 ,\I_5/plusOp__2_n_144 ,\I_5/plusOp__2_n_145 ,\I_5/plusOp__2_n_146 ,\I_5/plusOp__2_n_147 ,\I_5/plusOp__2_n_148 ,\I_5/plusOp__2_n_149 ,\I_5/plusOp__2_n_150 ,\I_5/plusOp__2_n_151 ,\I_5/plusOp__2_n_152 ,\I_5/plusOp__2_n_153 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__3_i_1 
       (.CI(\I_5/plusOp__3_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[2][10] ,\I_5/sr_reg_n_0_[2][9] ,\I_5/sr_reg_n_0_[2][8] }),
        .O({\I_5/plusOp__3_i_1_n_4 ,\I_5/plusOp__3_i_1_n_5 ,\I_5/plusOp__3_i_1_n_6 ,\I_5/plusOp__3_i_1_n_7 }),
        .S({\I_5/plusOp__3_i_4_n_0 ,\I_5/plusOp__3_i_5_n_0 ,\I_5/plusOp__3_i_6_n_0 ,\I_5/plusOp__3_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_10 
       (.I0(\I_5/sr_reg_n_0_[2][5] ),
        .I1(\I_5/sr_reg_n_0_[11][5] ),
        .O(\I_5/plusOp__3_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_11 
       (.I0(\I_5/sr_reg_n_0_[2][4] ),
        .I1(\I_5/sr_reg_n_0_[11][4] ),
        .O(\I_5/plusOp__3_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_12 
       (.I0(\I_5/sr_reg_n_0_[2][3] ),
        .I1(\I_5/sr_reg_n_0_[11][3] ),
        .O(\I_5/plusOp__3_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_13 
       (.I0(\I_5/sr_reg_n_0_[2][2] ),
        .I1(\I_5/sr_reg_n_0_[11][2] ),
        .O(\I_5/plusOp__3_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_14 
       (.I0(\I_5/sr_reg_n_0_[2][1] ),
        .I1(\I_5/sr_reg_n_0_[11][1] ),
        .O(\I_5/plusOp__3_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_15 
       (.I0(\I_5/sr_reg_n_0_[2][0] ),
        .I1(\I_5/sr_reg_n_0_[11][0] ),
        .O(\I_5/plusOp__3_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__3_i_2 
       (.CI(\I_5/plusOp__3_i_3_n_0 ),
        .CO({\I_5/plusOp__3_i_2_n_0 ,\I_5/plusOp__3_i_2_n_1 ,\I_5/plusOp__3_i_2_n_2 ,\I_5/plusOp__3_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[2][7] ,\I_5/sr_reg_n_0_[2][6] ,\I_5/sr_reg_n_0_[2][5] ,\I_5/sr_reg_n_0_[2][4] }),
        .O({\I_5/plusOp__3_i_2_n_4 ,\I_5/plusOp__3_i_2_n_5 ,\I_5/plusOp__3_i_2_n_6 ,\I_5/plusOp__3_i_2_n_7 }),
        .S({\I_5/plusOp__3_i_8_n_0 ,\I_5/plusOp__3_i_9_n_0 ,\I_5/plusOp__3_i_10_n_0 ,\I_5/plusOp__3_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp__3_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp__3_i_3_n_0 ,\I_5/plusOp__3_i_3_n_1 ,\I_5/plusOp__3_i_3_n_2 ,\I_5/plusOp__3_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[2][3] ,\I_5/sr_reg_n_0_[2][2] ,\I_5/sr_reg_n_0_[2][1] ,\I_5/sr_reg_n_0_[2][0] }),
        .O({\I_5/plusOp__3_i_3_n_4 ,\I_5/plusOp__3_i_3_n_5 ,\I_5/plusOp__3_i_3_n_6 ,\I_5/plusOp__3_i_3_n_7 }),
        .S({\I_5/plusOp__3_i_12_n_0 ,\I_5/plusOp__3_i_13_n_0 ,\I_5/plusOp__3_i_14_n_0 ,\I_5/plusOp__3_i_15_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_4 
       (.I0(\I_5/sr_reg_n_0_[2][11] ),
        .I1(\I_5/sr_reg_n_0_[11][11] ),
        .O(\I_5/plusOp__3_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_5 
       (.I0(\I_5/sr_reg_n_0_[2][10] ),
        .I1(\I_5/sr_reg_n_0_[11][10] ),
        .O(\I_5/plusOp__3_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_6 
       (.I0(\I_5/sr_reg_n_0_[2][9] ),
        .I1(\I_5/sr_reg_n_0_[11][9] ),
        .O(\I_5/plusOp__3_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_7 
       (.I0(\I_5/sr_reg_n_0_[2][8] ),
        .I1(\I_5/sr_reg_n_0_[11][8] ),
        .O(\I_5/plusOp__3_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_8 
       (.I0(\I_5/sr_reg_n_0_[2][7] ),
        .I1(\I_5/sr_reg_n_0_[11][7] ),
        .O(\I_5/plusOp__3_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \I_5/plusOp__3_i_9 
       (.I0(\I_5/sr_reg_n_0_[2][6] ),
        .I1(\I_5/sr_reg_n_0_[11][6] ),
        .O(\I_5/plusOp__3_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__3_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp_inferred__3_carry_n_0 ,\I_5/plusOp_inferred__3_carry_n_1 ,\I_5/plusOp_inferred__3_carry_n_2 ,\I_5/plusOp_inferred__3_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[14][3] ,\I_5/sr_reg_n_0_[14][2] ,\I_5/sr_reg_n_0_[14][1] ,\I_5/sr_reg_n_0_[14][0] }),
        .O({\I_5/plusOp_inferred__3_carry_n_4 ,\I_5/plusOp_inferred__3_carry_n_5 ,\I_5/plusOp_inferred__3_carry_n_6 ,\I_5/plusOp_inferred__3_carry_n_7 }),
        .S({plusOp_inferred__3_carry_i_1_n_0,plusOp_inferred__3_carry_i_2_n_0,plusOp_inferred__3_carry_i_3_n_0,plusOp_inferred__3_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__3_carry__0 
       (.CI(\I_5/plusOp_inferred__3_carry_n_0 ),
        .CO({\I_5/plusOp_inferred__3_carry__0_n_0 ,\I_5/plusOp_inferred__3_carry__0_n_1 ,\I_5/plusOp_inferred__3_carry__0_n_2 ,\I_5/plusOp_inferred__3_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[14][7] ,\I_5/sr_reg_n_0_[14][6] ,\I_5/sr_reg_n_0_[14][5] ,\I_5/sr_reg_n_0_[14][4] }),
        .O({\I_5/plusOp_inferred__3_carry__0_n_4 ,\I_5/plusOp_inferred__3_carry__0_n_5 ,\I_5/plusOp_inferred__3_carry__0_n_6 ,\I_5/plusOp_inferred__3_carry__0_n_7 }),
        .S({plusOp_inferred__3_carry__0_i_1_n_0,plusOp_inferred__3_carry__0_i_2_n_0,plusOp_inferred__3_carry__0_i_3_n_0,plusOp_inferred__3_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__3_carry__1 
       (.CI(\I_5/plusOp_inferred__3_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[14][10] ,\I_5/sr_reg_n_0_[14][9] ,\I_5/sr_reg_n_0_[14][8] }),
        .O({\I_5/plusOp_inferred__3_carry__1_n_4 ,\I_5/plusOp_inferred__3_carry__1_n_5 ,\I_5/plusOp_inferred__3_carry__1_n_6 ,\I_5/plusOp_inferred__3_carry__1_n_7 }),
        .S({plusOp_inferred__3_carry__1_i_1_n_0,plusOp_inferred__3_carry__1_i_2_n_0,plusOp_inferred__3_carry__1_i_3_n_0,plusOp_inferred__3_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__5_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp_inferred__5_carry_n_0 ,\I_5/plusOp_inferred__5_carry_n_1 ,\I_5/plusOp_inferred__5_carry_n_2 ,\I_5/plusOp_inferred__5_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[1][3] ,\I_5/sr_reg_n_0_[1][2] ,\I_5/sr_reg_n_0_[1][1] ,\I_5/sr_reg_n_0_[1][0] }),
        .O(\I_5/multOp__0 [3:0]),
        .S({plusOp_inferred__5_carry_i_1_n_0,plusOp_inferred__5_carry_i_2_n_0,plusOp_inferred__5_carry_i_3_n_0,plusOp_inferred__5_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__5_carry__0 
       (.CI(\I_5/plusOp_inferred__5_carry_n_0 ),
        .CO({\I_5/plusOp_inferred__5_carry__0_n_0 ,\I_5/plusOp_inferred__5_carry__0_n_1 ,\I_5/plusOp_inferred__5_carry__0_n_2 ,\I_5/plusOp_inferred__5_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[1][7] ,\I_5/sr_reg_n_0_[1][6] ,\I_5/sr_reg_n_0_[1][5] ,\I_5/sr_reg_n_0_[1][4] }),
        .O(\I_5/multOp__0 [7:4]),
        .S({plusOp_inferred__5_carry__0_i_1_n_0,plusOp_inferred__5_carry__0_i_2_n_0,plusOp_inferred__5_carry__0_i_3_n_0,plusOp_inferred__5_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__5_carry__1 
       (.CI(\I_5/plusOp_inferred__5_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[1][10] ,\I_5/sr_reg_n_0_[1][9] ,\I_5/sr_reg_n_0_[1][8] }),
        .O(\I_5/multOp__0 [11:8]),
        .S({plusOp_inferred__5_carry__1_i_1_n_0,plusOp_inferred__5_carry__1_i_2_n_0,plusOp_inferred__5_carry__1_i_3_n_0,plusOp_inferred__5_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__6_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp_inferred__6_carry_n_0 ,\I_5/plusOp_inferred__6_carry_n_1 ,\I_5/plusOp_inferred__6_carry_n_2 ,\I_5/plusOp_inferred__6_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[0][3] ,\I_5/sr_reg_n_0_[0][2] ,\I_5/sr_reg_n_0_[0][1] ,\I_5/sr_reg_n_0_ }),
        .O({\I_5/plusOp_inferred__6_carry_n_4 ,\I_5/plusOp_inferred__6_carry_n_5 ,\I_5/plusOp_inferred__6_carry_n_6 ,\I_5/plusOp_inferred__6_carry_n_7 }),
        .S({plusOp_inferred__6_carry_i_1_n_0,plusOp_inferred__6_carry_i_2_n_0,plusOp_inferred__6_carry_i_3_n_0,plusOp_inferred__6_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__6_carry__0 
       (.CI(\I_5/plusOp_inferred__6_carry_n_0 ),
        .CO({\I_5/plusOp_inferred__6_carry__0_n_0 ,\I_5/plusOp_inferred__6_carry__0_n_1 ,\I_5/plusOp_inferred__6_carry__0_n_2 ,\I_5/plusOp_inferred__6_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/sr_reg_n_0_[0][7] ,\I_5/sr_reg_n_0_[0][6] ,\I_5/sr_reg_n_0_[0][5] ,\I_5/sr_reg_n_0_[0][4] }),
        .O({\I_5/plusOp_inferred__6_carry__0_n_4 ,\I_5/plusOp_inferred__6_carry__0_n_5 ,\I_5/plusOp_inferred__6_carry__0_n_6 ,\I_5/plusOp_inferred__6_carry__0_n_7 }),
        .S({plusOp_inferred__6_carry__0_i_1_n_0,plusOp_inferred__6_carry__0_i_2_n_0,plusOp_inferred__6_carry__0_i_3_n_0,plusOp_inferred__6_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__6_carry__1 
       (.CI(\I_5/plusOp_inferred__6_carry__0_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_5/sr_reg_n_0_[0][10] ,\I_5/sr_reg_n_0_[0][9] ,\I_5/sr_reg_n_0_[0][8] }),
        .O({\I_5/plusOp_inferred__6_carry__1_n_4 ,\I_5/plusOp_inferred__6_carry__1_n_5 ,\I_5/plusOp_inferred__6_carry__1_n_6 ,\I_5/plusOp_inferred__6_carry__1_n_7 }),
        .S({plusOp_inferred__6_carry__1_i_1_n_0,plusOp_inferred__6_carry__1_i_2_n_0,plusOp_inferred__6_carry__1_i_3_n_0,plusOp_inferred__6_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp_inferred__7__62_carry_n_0 ,\I_5/plusOp_inferred__7__62_carry_n_1 ,\I_5/plusOp_inferred__7__62_carry_n_2 ,\I_5/plusOp_inferred__7__62_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/multOp__39_carry_n_7 ,\I_5/multOp_carry_n_5 ,\I_5/multOp_carry_n_6 ,\I_5/multOp_carry_n_7 }),
        .S({plusOp_inferred__7__62_carry_i_1_n_0,plusOp_inferred__7__62_carry_i_2_n_0,plusOp_inferred__7__62_carry_i_3_n_0,plusOp_inferred__7__62_carry_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry__0 
       (.CI(\I_5/plusOp_inferred__7__62_carry_n_0 ),
        .CO({\I_5/plusOp_inferred__7__62_carry__0_n_0 ,\I_5/plusOp_inferred__7__62_carry__0_n_1 ,\I_5/plusOp_inferred__7__62_carry__0_n_2 ,\I_5/plusOp_inferred__7__62_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/multOp__39_carry__0_n_7 ,\I_5/multOp__39_carry_n_4 ,\I_5/multOp__39_carry_n_5 ,\I_5/multOp__39_carry_n_6 }),
        .S({plusOp_inferred__7__62_carry__0_i_1_n_0,plusOp_inferred__7__62_carry__0_i_2_n_0,plusOp_inferred__7__62_carry__0_i_3_n_0,plusOp_inferred__7__62_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry__1 
       (.CI(\I_5/plusOp_inferred__7__62_carry__0_n_0 ),
        .CO({\I_5/plusOp_inferred__7__62_carry__1_n_0 ,\I_5/plusOp_inferred__7__62_carry__1_n_1 ,\I_5/plusOp_inferred__7__62_carry__1_n_2 ,\I_5/plusOp_inferred__7__62_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/multOp__39_carry__1_n_7 ,\I_5/multOp__39_carry__0_n_4 ,\I_5/multOp__39_carry__0_n_5 ,\I_5/multOp__39_carry__0_n_6 }),
        .O({\I_5/plusOp_inferred__7__62_carry__1_n_4 ,\I_5/plusOp_inferred__7__62_carry__1_n_5 ,\I_5/plusOp_inferred__7__62_carry__1_n_6 ,\I_5/plusOp_inferred__7__62_carry__1_n_7 }),
        .S({plusOp_inferred__7__62_carry__1_i_1_n_0,plusOp_inferred__7__62_carry__1_i_2_n_0,plusOp_inferred__7__62_carry__1_i_3_n_0,plusOp_inferred__7__62_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry__2 
       (.CI(\I_5/plusOp_inferred__7__62_carry__1_n_0 ),
        .CO({\I_5/plusOp_inferred__7__62_carry__2_n_0 ,\I_5/plusOp_inferred__7__62_carry__2_n_1 ,\I_5/plusOp_inferred__7__62_carry__2_n_2 ,\I_5/plusOp_inferred__7__62_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({plusOp_inferred__7__62_carry__2_i_1_n_0,\I_5/multOp__39_carry__1_n_4 ,\I_5/multOp__39_carry__1_n_5 ,\I_5/multOp__39_carry__1_n_6 }),
        .O({\I_5/plusOp_inferred__7__62_carry__2_n_4 ,\I_5/plusOp_inferred__7__62_carry__2_n_5 ,\I_5/plusOp_inferred__7__62_carry__2_n_6 ,\I_5/plusOp_inferred__7__62_carry__2_n_7 }),
        .S({plusOp_inferred__7__62_carry__2_i_2_n_0,plusOp_inferred__7__62_carry__2_i_3_n_0,plusOp_inferred__7__62_carry__2_i_4_n_0,plusOp_inferred__7__62_carry__2_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry__3 
       (.CI(\I_5/plusOp_inferred__7__62_carry__2_n_0 ),
        .CO({\I_5/plusOp_inferred__7__62_carry__3_n_0 ,\I_5/plusOp_inferred__7__62_carry__3_n_1 ,\I_5/plusOp_inferred__7__62_carry__3_n_2 ,\I_5/plusOp_inferred__7__62_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(C[18:15]),
        .O({\I_5/plusOp_inferred__7__62_carry__3_n_4 ,\I_5/plusOp_inferred__7__62_carry__3_n_5 ,\I_5/plusOp_inferred__7__62_carry__3_n_6 ,\I_5/plusOp_inferred__7__62_carry__3_n_7 }),
        .S({plusOp_inferred__7__62_carry__3_i_1_n_0,plusOp_inferred__7__62_carry__3_i_2_n_0,plusOp_inferred__7__62_carry__3_i_3_n_0,plusOp_inferred__7__62_carry__3_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7__62_carry__4 
       (.CI(\I_5/plusOp_inferred__7__62_carry__3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,C[20:19]}),
        .O({\I_5/plusOp_inferred__7__62_carry__4_n_4 ,\I_5/plusOp_inferred__7__62_carry__4_n_5 ,\I_5/plusOp_inferred__7__62_carry__4_n_6 ,\I_5/plusOp_inferred__7__62_carry__4_n_7 }),
        .S({\<const0>__0__0 ,plusOp_inferred__7__62_carry__4_i_1_n_0,plusOp_inferred__7__62_carry__4_i_2_n_0,plusOp_inferred__7__62_carry__4_i_3_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry 
       (.CI(\<const0>__0__0 ),
        .CO({\I_5/plusOp_inferred__7_carry_n_0 ,\I_5/plusOp_inferred__7_carry_n_1 ,\I_5/plusOp_inferred__7_carry_n_2 ,\I_5/plusOp_inferred__7_carry_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/multOp__0 [2:0],\<const0>__0__0 }),
        .O(C[4:1]),
        .S({plusOp_inferred__7_carry_i_1_n_0,plusOp_inferred__7_carry_i_2_n_0,plusOp_inferred__7_carry_i_3_n_0,\I_5/plusOp__3_n_104 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry__0 
       (.CI(\I_5/plusOp_inferred__7_carry_n_0 ),
        .CO({\I_5/plusOp_inferred__7_carry__0_n_0 ,\I_5/plusOp_inferred__7_carry__0_n_1 ,\I_5/plusOp_inferred__7_carry__0_n_2 ,\I_5/plusOp_inferred__7_carry__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_5/multOp__0 [6:3]),
        .O(C[8:5]),
        .S({plusOp_inferred__7_carry__0_i_1_n_0,plusOp_inferred__7_carry__0_i_2_n_0,plusOp_inferred__7_carry__0_i_3_n_0,plusOp_inferred__7_carry__0_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry__1 
       (.CI(\I_5/plusOp_inferred__7_carry__0_n_0 ),
        .CO({\I_5/plusOp_inferred__7_carry__1_n_0 ,\I_5/plusOp_inferred__7_carry__1_n_1 ,\I_5/plusOp_inferred__7_carry__1_n_2 ,\I_5/plusOp_inferred__7_carry__1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_5/multOp__0 [10:7]),
        .O(C[12:9]),
        .S({plusOp_inferred__7_carry__1_i_1_n_0,plusOp_inferred__7_carry__1_i_2_n_0,plusOp_inferred__7_carry__1_i_3_n_0,plusOp_inferred__7_carry__1_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry__2 
       (.CI(\I_5/plusOp_inferred__7_carry__1_n_0 ),
        .CO({\I_5/plusOp_inferred__7_carry__2_n_0 ,\I_5/plusOp_inferred__7_carry__2_n_1 ,\I_5/plusOp_inferred__7_carry__2_n_2 ,\I_5/plusOp_inferred__7_carry__2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/plusOp__3_n_90 ,\I_5/plusOp__3_n_91 ,\I_5/plusOp__3_n_92 ,plusOp_inferred__7_carry__2_i_1_n_0}),
        .O(C[16:13]),
        .S({plusOp_inferred__7_carry__2_i_2_n_0,plusOp_inferred__7_carry__2_i_3_n_0,plusOp_inferred__7_carry__2_i_4_n_0,plusOp_inferred__7_carry__2_i_5_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry__3 
       (.CI(\I_5/plusOp_inferred__7_carry__2_n_0 ),
        .CO({\I_5/plusOp_inferred__7_carry__3_n_0 ,\I_5/plusOp_inferred__7_carry__3_n_1 ,\I_5/plusOp_inferred__7_carry__3_n_2 ,\I_5/plusOp_inferred__7_carry__3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_5/plusOp__3_n_86 ,\I_5/plusOp__3_n_87 ,\I_5/plusOp__3_n_88 ,\I_5/plusOp__3_n_89 }),
        .O(C[20:17]),
        .S({plusOp_inferred__7_carry__3_i_1_n_0,plusOp_inferred__7_carry__3_i_2_n_0,plusOp_inferred__7_carry__3_i_3_n_0,plusOp_inferred__7_carry__3_i_4_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \I_5/plusOp_inferred__7_carry__4 
       (.CI(\I_5/plusOp_inferred__7_carry__3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_5/plusOp__3_n_85 }),
        .O({\I_5/plusOp_inferred__7_carry__4_n_4 ,\I_5/plusOp_inferred__7_carry__4_n_5 ,C[22:21]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,plusOp_inferred__7_carry__4_i_1_n_0,plusOp_inferred__7_carry__4_i_2_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[0]),
        .Q(\I_5/sr_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(pre_yuv_v[10]),
        .Q(\I_5/sr_reg_n_0_[0][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(pre_yuv_v[11]),
        .Q(\I_5/sr_reg_n_0_[0][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[1]),
        .Q(\I_5/sr_reg_n_0_[0][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[2]),
        .Q(\I_5/sr_reg_n_0_[0][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[3]),
        .Q(\I_5/sr_reg_n_0_[0][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[4]),
        .Q(\I_5/sr_reg_n_0_[0][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[5]),
        .Q(\I_5/sr_reg_n_0_[0][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[6]),
        .Q(\I_5/sr_reg_n_0_[0][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(pre_yuv_v[7]),
        .Q(\I_5/sr_reg_n_0_[0][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(pre_yuv_v[8]),
        .Q(\I_5/sr_reg_n_0_[0][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[0][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(pre_yuv_v[9]),
        .Q(\I_5/sr_reg_n_0_[0][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][0] ),
        .Q(\I_5/sr_reg_n_0_[10][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][10] ),
        .Q(\I_5/sr_reg_n_0_[10][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][11] ),
        .Q(\I_5/sr_reg_n_0_[10][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][1] ),
        .Q(\I_5/sr_reg_n_0_[10][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][2] ),
        .Q(\I_5/sr_reg_n_0_[10][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][3] ),
        .Q(\I_5/sr_reg_n_0_[10][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[9][4] ),
        .Q(\I_5/sr_reg_n_0_[10][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[9][5] ),
        .Q(\I_5/sr_reg_n_0_[10][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[9][6] ),
        .Q(\I_5/sr_reg_n_0_[10][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[9][7] ),
        .Q(\I_5/sr_reg_n_0_[10][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][8] ),
        .Q(\I_5/sr_reg_n_0_[10][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[10][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[9][9] ),
        .Q(\I_5/sr_reg_n_0_[10][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][0] ),
        .Q(\I_5/sr_reg_n_0_[11][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[10][10] ),
        .Q(\I_5/sr_reg_n_0_[11][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[10][11] ),
        .Q(\I_5/sr_reg_n_0_[11][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][1] ),
        .Q(\I_5/sr_reg_n_0_[11][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][2] ),
        .Q(\I_5/sr_reg_n_0_[11][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][3] ),
        .Q(\I_5/sr_reg_n_0_[11][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][4] ),
        .Q(\I_5/sr_reg_n_0_[11][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][5] ),
        .Q(\I_5/sr_reg_n_0_[11][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][6] ),
        .Q(\I_5/sr_reg_n_0_[11][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[10][7] ),
        .Q(\I_5/sr_reg_n_0_[11][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[10][8] ),
        .Q(\I_5/sr_reg_n_0_[11][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[11][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[10][9] ),
        .Q(\I_5/sr_reg_n_0_[11][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][0] ),
        .Q(\I_5/sr_reg_n_0_[12][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][10] ),
        .Q(\I_5/sr_reg_n_0_[12][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][11] ),
        .Q(\I_5/sr_reg_n_0_[12][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][1] ),
        .Q(\I_5/sr_reg_n_0_[12][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][2] ),
        .Q(\I_5/sr_reg_n_0_[12][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][3] ),
        .Q(\I_5/sr_reg_n_0_[12][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][4] ),
        .Q(\I_5/sr_reg_n_0_[12][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][5] ),
        .Q(\I_5/sr_reg_n_0_[12][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][6] ),
        .Q(\I_5/sr_reg_n_0_[12][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][7] ),
        .Q(\I_5/sr_reg_n_0_[12][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][8] ),
        .Q(\I_5/sr_reg_n_0_[12][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[12][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[11][9] ),
        .Q(\I_5/sr_reg_n_0_[12][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][0] ),
        .Q(\I_5/sr_reg_n_0_[13][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[12][10] ),
        .Q(\I_5/sr_reg_n_0_[13][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[12][11] ),
        .Q(\I_5/sr_reg_n_0_[13][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][1] ),
        .Q(\I_5/sr_reg_n_0_[13][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][2] ),
        .Q(\I_5/sr_reg_n_0_[13][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][3] ),
        .Q(\I_5/sr_reg_n_0_[13][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][4] ),
        .Q(\I_5/sr_reg_n_0_[13][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][5] ),
        .Q(\I_5/sr_reg_n_0_[13][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][6] ),
        .Q(\I_5/sr_reg_n_0_[13][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[12][7] ),
        .Q(\I_5/sr_reg_n_0_[13][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[12][8] ),
        .Q(\I_5/sr_reg_n_0_[13][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[13][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[12][9] ),
        .Q(\I_5/sr_reg_n_0_[13][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][0] ),
        .Q(\I_5/sr_reg_n_0_[14][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][10] ),
        .Q(\I_5/sr_reg_n_0_[14][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][11] ),
        .Q(\I_5/sr_reg_n_0_[14][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][1] ),
        .Q(\I_5/sr_reg_n_0_[14][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][2] ),
        .Q(\I_5/sr_reg_n_0_[14][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][3] ),
        .Q(\I_5/sr_reg_n_0_[14][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][4] ),
        .Q(\I_5/sr_reg_n_0_[14][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][5] ),
        .Q(\I_5/sr_reg_n_0_[14][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][6] ),
        .Q(\I_5/sr_reg_n_0_[14][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][7] ),
        .Q(\I_5/sr_reg_n_0_[14][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][8] ),
        .Q(\I_5/sr_reg_n_0_[14][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[14][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[13][9] ),
        .Q(\I_5/sr_reg_n_0_[14][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_ ),
        .Q(\I_5/sr_reg_n_0_[1][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[0][10] ),
        .Q(\I_5/sr_reg_n_0_[1][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[0][11] ),
        .Q(\I_5/sr_reg_n_0_[1][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][1] ),
        .Q(\I_5/sr_reg_n_0_[1][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][2] ),
        .Q(\I_5/sr_reg_n_0_[1][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][3] ),
        .Q(\I_5/sr_reg_n_0_[1][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][4] ),
        .Q(\I_5/sr_reg_n_0_[1][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][5] ),
        .Q(\I_5/sr_reg_n_0_[1][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][6] ),
        .Q(\I_5/sr_reg_n_0_[1][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\I_5/sr_reg_n_0_[0][7] ),
        .Q(\I_5/sr_reg_n_0_[1][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[0][8] ),
        .Q(\I_5/sr_reg_n_0_[1][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[1][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(en_bild_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[0][9] ),
        .Q(\I_5/sr_reg_n_0_[1][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][0] ),
        .Q(\I_5/sr_reg_n_0_[2][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][10] ),
        .Q(\I_5/sr_reg_n_0_[2][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][11] ),
        .Q(\I_5/sr_reg_n_0_[2][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][1] ),
        .Q(\I_5/sr_reg_n_0_[2][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][2] ),
        .Q(\I_5/sr_reg_n_0_[2][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][3] ),
        .Q(\I_5/sr_reg_n_0_[2][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[1][4] ),
        .Q(\I_5/sr_reg_n_0_[2][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[1][5] ),
        .Q(\I_5/sr_reg_n_0_[2][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[1][6] ),
        .Q(\I_5/sr_reg_n_0_[2][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[1][7] ),
        .Q(\I_5/sr_reg_n_0_[2][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][8] ),
        .Q(\I_5/sr_reg_n_0_[2][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[2][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[1][9] ),
        .Q(\I_5/sr_reg_n_0_[2][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][0] ),
        .Q(\I_5/sr_reg_n_0_[3][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][10] ),
        .Q(\I_5/sr_reg_n_0_[3][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][11] ),
        .Q(\I_5/sr_reg_n_0_[3][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][1] ),
        .Q(\I_5/sr_reg_n_0_[3][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][2] ),
        .Q(\I_5/sr_reg_n_0_[3][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][3] ),
        .Q(\I_5/sr_reg_n_0_[3][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[2][4] ),
        .Q(\I_5/sr_reg_n_0_[3][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[2][5] ),
        .Q(\I_5/sr_reg_n_0_[3][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[2][6] ),
        .Q(\I_5/sr_reg_n_0_[3][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[2][7] ),
        .Q(\I_5/sr_reg_n_0_[3][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][8] ),
        .Q(\I_5/sr_reg_n_0_[3][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[3][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[2][9] ),
        .Q(\I_5/sr_reg_n_0_[3][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][0] ),
        .Q(\I_5/sr_reg_n_0_[4][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][10] ),
        .Q(\I_5/sr_reg_n_0_[4][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][11] ),
        .Q(\I_5/sr_reg_n_0_[4][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][1] ),
        .Q(\I_5/sr_reg_n_0_[4][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][2] ),
        .Q(\I_5/sr_reg_n_0_[4][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][3] ),
        .Q(\I_5/sr_reg_n_0_[4][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[3][4] ),
        .Q(\I_5/sr_reg_n_0_[4][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[3][5] ),
        .Q(\I_5/sr_reg_n_0_[4][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[3][6] ),
        .Q(\I_5/sr_reg_n_0_[4][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[3][7] ),
        .Q(\I_5/sr_reg_n_0_[4][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][8] ),
        .Q(\I_5/sr_reg_n_0_[4][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[4][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[3][9] ),
        .Q(\I_5/sr_reg_n_0_[4][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][0] ),
        .Q(\I_5/sr_reg_n_0_[5][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][10] ),
        .Q(\I_5/sr_reg_n_0_[5][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][11] ),
        .Q(\I_5/sr_reg_n_0_[5][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][1] ),
        .Q(\I_5/sr_reg_n_0_[5][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][2] ),
        .Q(\I_5/sr_reg_n_0_[5][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][3] ),
        .Q(\I_5/sr_reg_n_0_[5][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[4][4] ),
        .Q(\I_5/sr_reg_n_0_[5][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[4][5] ),
        .Q(\I_5/sr_reg_n_0_[5][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[4][6] ),
        .Q(\I_5/sr_reg_n_0_[5][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[4][7] ),
        .Q(\I_5/sr_reg_n_0_[5][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][8] ),
        .Q(\I_5/sr_reg_n_0_[5][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[5][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[4][9] ),
        .Q(\I_5/sr_reg_n_0_[5][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][0] ),
        .Q(\I_5/sr_reg_n_0_[6][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][10] ),
        .Q(\I_5/sr_reg_n_0_[6][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][11] ),
        .Q(\I_5/sr_reg_n_0_[6][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][1] ),
        .Q(\I_5/sr_reg_n_0_[6][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][2] ),
        .Q(\I_5/sr_reg_n_0_[6][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][3] ),
        .Q(\I_5/sr_reg_n_0_[6][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[5][4] ),
        .Q(\I_5/sr_reg_n_0_[6][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[5][5] ),
        .Q(\I_5/sr_reg_n_0_[6][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[5][6] ),
        .Q(\I_5/sr_reg_n_0_[6][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[5][7] ),
        .Q(\I_5/sr_reg_n_0_[6][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][8] ),
        .Q(\I_5/sr_reg_n_0_[6][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[6][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[5][9] ),
        .Q(\I_5/sr_reg_n_0_[6][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][0] ),
        .Q(\I_5/sr_reg_n_0_[7][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][10] ),
        .Q(\I_5/sr_reg_n_0_[7][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][11] ),
        .Q(\I_5/sr_reg_n_0_[7][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][1] ),
        .Q(\I_5/sr_reg_n_0_[7][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][2] ),
        .Q(\I_5/sr_reg_n_0_[7][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][3] ),
        .Q(\I_5/sr_reg_n_0_[7][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[6][4] ),
        .Q(\I_5/sr_reg_n_0_[7][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[6][5] ),
        .Q(\I_5/sr_reg_n_0_[7][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[6][6] ),
        .Q(\I_5/sr_reg_n_0_[7][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[6][7] ),
        .Q(\I_5/sr_reg_n_0_[7][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][8] ),
        .Q(\I_5/sr_reg_n_0_[7][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[7][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[6][9] ),
        .Q(\I_5/sr_reg_n_0_[7][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][0] ),
        .Q(\I_5/sr_reg_n_0_[8][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][10] ),
        .Q(\I_5/sr_reg_n_0_[8][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][11] ),
        .Q(\I_5/sr_reg_n_0_[8][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][1] ),
        .Q(\I_5/sr_reg_n_0_[8][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][2] ),
        .Q(\I_5/sr_reg_n_0_[8][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][3] ),
        .Q(\I_5/sr_reg_n_0_[8][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[7][4] ),
        .Q(\I_5/sr_reg_n_0_[8][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[7][5] ),
        .Q(\I_5/sr_reg_n_0_[8][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[7][6] ),
        .Q(\I_5/sr_reg_n_0_[8][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[7][7] ),
        .Q(\I_5/sr_reg_n_0_[8][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][8] ),
        .Q(\I_5/sr_reg_n_0_[8][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[8][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[7][9] ),
        .Q(\I_5/sr_reg_n_0_[8][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][0] ),
        .Q(\I_5/sr_reg_n_0_[9][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][10] ),
        .Q(\I_5/sr_reg_n_0_[9][10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][11] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][11] ),
        .Q(\I_5/sr_reg_n_0_[9][11] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][1] ),
        .Q(\I_5/sr_reg_n_0_[9][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][2] ),
        .Q(\I_5/sr_reg_n_0_[9][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][3] ),
        .Q(\I_5/sr_reg_n_0_[9][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[8][4] ),
        .Q(\I_5/sr_reg_n_0_[9][4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[8][5] ),
        .Q(\I_5/sr_reg_n_0_[9][5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[8][6] ),
        .Q(\I_5/sr_reg_n_0_[9][6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(\sr[2][7]_i_1_n_0 ),
        .D(\I_5/sr_reg_n_0_[8][7] ),
        .Q(\I_5/sr_reg_n_0_[9][7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][8] ),
        .Q(\I_5/sr_reg_n_0_[9][8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_5/sr_reg[9][9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_5/sr_reg_n_0_[8][9] ),
        .Q(\I_5/sr_reg_n_0_[9][9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[0] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__9_n_0 ),
        .Q(\I_6/output_reg_n_0_ ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[10] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate_n_0 ),
        .Q(\I_6/output_reg_n_0_[10] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[1] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__8_n_0 ),
        .Q(\I_6/output_reg_n_0_[1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[2] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__7_n_0 ),
        .Q(\I_6/output_reg_n_0_[2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[3] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__6_n_0 ),
        .Q(\I_6/output_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[4] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__5_n_0 ),
        .Q(\I_6/output_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[5] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__4_n_0 ),
        .Q(\I_6/output_reg_n_0_[5] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[6] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__3_n_0 ),
        .Q(\I_6/output_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[7] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__2_n_0 ),
        .Q(\I_6/output_reg_n_0_[7] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[8] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__1_n_0 ),
        .Q(\I_6/output_reg_n_0_[8] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/output_reg[9] 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_gate__0_n_0 ),
        .Q(\I_6/output_reg_n_0_[9] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][0]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][0]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[0]),
        .Q(\I_6/sr_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][10]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][10]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[10]),
        .Q(\I_6/sr_reg[5][10]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][1]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][1]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[1]),
        .Q(\I_6/sr_reg[5][1]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][2]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][2]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[2]),
        .Q(\I_6/sr_reg[5][2]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][3]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][3]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[3]),
        .Q(\I_6/sr_reg[5][3]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][4]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][4]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[4]),
        .Q(\I_6/sr_reg[5][4]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][5]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][5]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[5]),
        .Q(\I_6/sr_reg[5][5]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][6]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][6]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[6]),
        .Q(\I_6/sr_reg[5][6]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][7]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][7]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[7]),
        .Q(\I_6/sr_reg[5][7]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][8]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][8]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[8]),
        .Q(\I_6/sr_reg[5][8]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "graphiti_0/\I_6/sr_reg[5] " *) 
  (* srl_name = "graphiti_0/\I_6/sr_reg[5][9]_srl7_I_6_sr_reg_c_4 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \I_6/sr_reg[5][9]_srl7_I_6_sr_reg_c_4 
       (.A0(\<const0>__0__0 ),
        .A1(\<const1>__0__0 ),
        .A2(\<const1>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk15M),
        .D(plusOp18[9]),
        .Q(\I_6/sr_reg[5][9]_srl7_I_6_sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][0]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg ),
        .Q(\I_6/sr_reg[6][0]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][10]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][10]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][10]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][1]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][1]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][1]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][2]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][2]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][2]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][3]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][3]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][3]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][4]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][4]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][4]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][5]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][5]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][5]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][6]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][6]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][6]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][7]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][7]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][7]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][8]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][8]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][8]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \I_6/sr_reg[6][9]_I_6_sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .D(\I_6/sr_reg[5][9]_srl7_I_6_sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg[6][9]_I_6_sr_reg_c_5_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_3/out_y_reg_c_n_0 ),
        .Q(\I_6/sr_reg_c_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_0 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_n_0 ),
        .Q(\I_6/sr_reg_c_0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_1 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_0_n_0 ),
        .Q(\I_6/sr_reg_c_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_2 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_1_n_0 ),
        .Q(\I_6/sr_reg_c_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_3 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_2_n_0 ),
        .Q(\I_6/sr_reg_c_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_4 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_3_n_0 ),
        .Q(\I_6/sr_reg_c_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \I_6/sr_reg_c_5 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(i_austastung_i_2_n_0),
        .D(\I_6/sr_reg_c_4_n_0 ),
        .Q(\I_6/sr_reg_c_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate 
       (.I0(\I_6/sr_reg[6][10]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__0 
       (.I0(\I_6/sr_reg[6][9]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__1 
       (.I0(\I_6/sr_reg[6][8]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__2 
       (.I0(\I_6/sr_reg[6][7]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__3 
       (.I0(\I_6/sr_reg[6][6]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__4 
       (.I0(\I_6/sr_reg[6][5]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__5 
       (.I0(\I_6/sr_reg[6][4]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__6 
       (.I0(\I_6/sr_reg[6][3]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__7 
       (.I0(\I_6/sr_reg[6][2]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__8 
       (.I0(\I_6/sr_reg[6][1]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \I_6/sr_reg_gate__9 
       (.I0(\I_6/sr_reg[6][0]_I_6_sr_reg_c_5_n_0 ),
        .I1(\I_6/sr_reg_c_5_n_0 ),
        .O(\I_6/sr_reg_gate__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_1
       (.P(VCC_2));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \abschnittu[1]_i_10 
       (.I0(\I_1/ctr_48_reg [56]),
        .O(\abschnittu[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \abschnittu[1]_i_5 
       (.I0(\I_1/ctr90_48_reg [60]),
        .O(\abschnittu[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \abschnittu[1]_i_6 
       (.I0(\I_1/ctr_48_reg [60]),
        .O(\abschnittu[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \abschnittu[1]_i_7 
       (.I0(\I_1/ctr_48_reg [59]),
        .O(\abschnittu[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \abschnittu_reg[1]_i_1 
       (.CI(adr_reg_i_16_n_0),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [60]}),
        .O({p_2_in,p_2_in__0[7:5]}),
        .S({\I_1/ctr90_48_reg [63:61],\abschnittu[1]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \abschnittu_reg[1]_i_1__0 
       (.CI(abschnittu_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [60]}),
        .O({p_3_in,p_3_in__0[7:5]}),
        .S({\I_1/ctr_48_reg [63:61],\abschnittu[1]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \abschnittu_reg[1]_i_2 
       (.CI(adr_reg_i_15_n_0),
        .CO(abschnittu_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr_48_reg [59],\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [56]}),
        .O(p_3_in__0[4:1]),
        .S({\abschnittu[1]_i_7_n_0 ,\I_1/ctr_48_reg [58:57],\abschnittu[1]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_100
       (.I0(\I_1/ctr90_48_reg [25]),
        .O(adr_reg_i_100_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_101
       (.I0(\I_1/ctr90_48_reg [24]),
        .O(adr_reg_i_101_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_102
       (.CI(adr_reg_i_112_n_0),
        .CO({adr_reg_i_102_n_0,adr_reg_i_102_n_1,adr_reg_i_102_n_2,adr_reg_i_102_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [16]}),
        .S({\I_1/ctr_48_reg [19:17],adr_reg_i_116_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_106
       (.I0(\I_1/ctr_48_reg [20]),
        .O(adr_reg_i_106_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_107
       (.CI(adr_reg_i_117_n_0),
        .CO({adr_reg_i_107_n_0,adr_reg_i_107_n_1,adr_reg_i_107_n_2,adr_reg_i_107_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [16]}),
        .S({\I_1/ctr90_48_reg [19:17],adr_reg_i_121_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_111
       (.I0(\I_1/ctr90_48_reg [20]),
        .O(adr_reg_i_111_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_112
       (.CI(adr_reg_i_122_n_0),
        .CO({adr_reg_i_112_n_0,adr_reg_i_112_n_1,adr_reg_i_112_n_2,adr_reg_i_112_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr_48_reg [14:12]}),
        .S({\I_1/ctr_48_reg [15],adr_reg_i_124_n_0,adr_reg_i_125_n_0,adr_reg_i_126_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_116
       (.I0(\I_1/ctr_48_reg [16]),
        .O(adr_reg_i_116_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_117
       (.CI(adr_reg_i_127_n_0),
        .CO({adr_reg_i_117_n_0,adr_reg_i_117_n_1,adr_reg_i_117_n_2,adr_reg_i_117_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr90_48_reg [14:12]}),
        .S({\I_1/ctr90_48_reg [15],adr_reg_i_129_n_0,adr_reg_i_130_n_0,adr_reg_i_131_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_121
       (.I0(\I_1/ctr90_48_reg [16]),
        .O(adr_reg_i_121_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_122
       (.CI(adr_reg_i_132_n_0),
        .CO({adr_reg_i_122_n_0,adr_reg_i_122_n_1,adr_reg_i_122_n_2,adr_reg_i_122_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr_48_reg [10],\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\I_1/ctr_48_reg [11],adr_reg_i_134_n_0,\I_1/ctr_48_reg [9:8]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_124
       (.I0(\I_1/ctr_48_reg [14]),
        .O(adr_reg_i_124_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_125
       (.I0(\I_1/ctr_48_reg [13]),
        .O(adr_reg_i_125_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_126
       (.I0(\I_1/ctr_48_reg [12]),
        .O(adr_reg_i_126_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_127
       (.CI(adr_reg_i_137_n_0),
        .CO({adr_reg_i_127_n_0,adr_reg_i_127_n_1,adr_reg_i_127_n_2,adr_reg_i_127_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr90_48_reg [10],\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\I_1/ctr90_48_reg [11],adr_reg_i_139_n_0,\I_1/ctr90_48_reg [9:8]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_129
       (.I0(\I_1/ctr90_48_reg [14]),
        .O(adr_reg_i_129_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_130
       (.I0(\I_1/ctr90_48_reg [13]),
        .O(adr_reg_i_130_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_131
       (.I0(\I_1/ctr90_48_reg [12]),
        .O(adr_reg_i_131_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_132
       (.CI(adr_reg_i_142_n_0),
        .CO({adr_reg_i_132_n_0,adr_reg_i_132_n_1,adr_reg_i_132_n_2,adr_reg_i_132_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_1/ctr_48_reg [7:4]),
        .S({adr_reg_i_143_n_0,adr_reg_i_144_n_0,adr_reg_i_145_n_0,adr_reg_i_146_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_134
       (.I0(\I_1/ctr_48_reg [10]),
        .O(adr_reg_i_134_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_137
       (.CI(adr_reg_i_147_n_0),
        .CO({adr_reg_i_137_n_0,adr_reg_i_137_n_1,adr_reg_i_137_n_2,adr_reg_i_137_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI(\I_1/ctr90_48_reg [7:4]),
        .S({adr_reg_i_148_n_0,adr_reg_i_149_n_0,adr_reg_i_150_n_0,adr_reg_i_151_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_139
       (.I0(\I_1/ctr90_48_reg [10]),
        .O(adr_reg_i_139_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_142
       (.CI(\<const0>__0__0 ),
        .CO({adr_reg_i_142_n_0,adr_reg_i_142_n_1,adr_reg_i_142_n_2,adr_reg_i_142_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [1],\<const0>__0__0 }),
        .S({\I_1/ctr_48_reg [3:2],adr_reg_i_154_n_0,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_143
       (.I0(\I_1/ctr_48_reg [7]),
        .O(adr_reg_i_143_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_144
       (.I0(\I_1/ctr_48_reg [6]),
        .O(adr_reg_i_144_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_145
       (.I0(\I_1/ctr_48_reg [5]),
        .O(adr_reg_i_145_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_146
       (.I0(\I_1/ctr_48_reg [4]),
        .O(adr_reg_i_146_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_147
       (.CI(\<const0>__0__0 ),
        .CO({adr_reg_i_147_n_0,adr_reg_i_147_n_1,adr_reg_i_147_n_2,adr_reg_i_147_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [1],\<const0>__0__0 }),
        .S({\I_1/ctr90_48_reg [3:2],adr_reg_i_157_n_0,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_148
       (.I0(\I_1/ctr90_48_reg [7]),
        .O(adr_reg_i_148_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_149
       (.I0(\I_1/ctr90_48_reg [6]),
        .O(adr_reg_i_149_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_15
       (.CI(adr_reg_i_18_n_0),
        .CO({adr_reg_i_15_n_0,adr_reg_i_15_n_1,adr_reg_i_15_n_2,adr_reg_i_15_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [53:52]}),
        .O({p_3_in__0[0],adr_reg_i_15_n_5,adr_reg_i_15_n_6,adr_reg_i_15_n_7}),
        .S({\I_1/ctr_48_reg [55:54],adr_reg_i_21_n_0,adr_reg_i_22_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_150
       (.I0(\I_1/ctr90_48_reg [5]),
        .O(adr_reg_i_150_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_151
       (.I0(\I_1/ctr90_48_reg [4]),
        .O(adr_reg_i_151_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_154
       (.I0(\I_1/ctr_48_reg [1]),
        .O(adr_reg_i_154_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_157
       (.I0(\I_1/ctr90_48_reg [1]),
        .O(adr_reg_i_157_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_16
       (.CI(adr_reg_i_17_n_0),
        .CO({adr_reg_i_16_n_0,adr_reg_i_16_n_1,adr_reg_i_16_n_2,adr_reg_i_16_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr90_48_reg [59],\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [56]}),
        .O(p_2_in__0[4:1]),
        .S({adr_reg_i_23_n_0,\I_1/ctr90_48_reg [58:57],adr_reg_i_26_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_17
       (.CI(adr_reg_i_27_n_0),
        .CO({adr_reg_i_17_n_0,adr_reg_i_17_n_1,adr_reg_i_17_n_2,adr_reg_i_17_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [53:52]}),
        .O({p_2_in__0[0],adr_reg_i_17_n_5,adr_reg_i_17_n_6,adr_reg_i_17_n_7}),
        .S({\I_1/ctr90_48_reg [55:54],adr_reg_i_30_n_0,adr_reg_i_31_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_18
       (.CI(adr_reg_i_32_n_0),
        .CO({adr_reg_i_18_n_0,adr_reg_i_18_n_1,adr_reg_i_18_n_2,adr_reg_i_18_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr_48_reg [51],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({adr_reg_i_33_n_0,\I_1/ctr_48_reg [50:48]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_21
       (.I0(\I_1/ctr_48_reg [53]),
        .O(adr_reg_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_22
       (.I0(\I_1/ctr_48_reg [52]),
        .O(adr_reg_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_23
       (.I0(\I_1/ctr90_48_reg [59]),
        .O(adr_reg_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_26
       (.I0(\I_1/ctr90_48_reg [56]),
        .O(adr_reg_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_27
       (.CI(adr_reg_i_37_n_0),
        .CO({adr_reg_i_27_n_0,adr_reg_i_27_n_1,adr_reg_i_27_n_2,adr_reg_i_27_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr90_48_reg [51],\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({adr_reg_i_38_n_0,\I_1/ctr90_48_reg [50:48]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_30
       (.I0(\I_1/ctr90_48_reg [53]),
        .O(adr_reg_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_31
       (.I0(\I_1/ctr90_48_reg [52]),
        .O(adr_reg_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_32
       (.CI(adr_reg_i_42_n_0),
        .CO({adr_reg_i_32_n_0,adr_reg_i_32_n_1,adr_reg_i_32_n_2,adr_reg_i_32_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr_48_reg [47:45],\<const0>__0__0 }),
        .S({adr_reg_i_43_n_0,adr_reg_i_44_n_0,adr_reg_i_45_n_0,\I_1/ctr_48_reg [44]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_33
       (.I0(\I_1/ctr_48_reg [51]),
        .O(adr_reg_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_37
       (.CI(adr_reg_i_47_n_0),
        .CO({adr_reg_i_37_n_0,adr_reg_i_37_n_1,adr_reg_i_37_n_2,adr_reg_i_37_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr90_48_reg [47:45],\<const0>__0__0 }),
        .S({adr_reg_i_48_n_0,adr_reg_i_49_n_0,adr_reg_i_50_n_0,\I_1/ctr90_48_reg [44]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_38
       (.I0(\I_1/ctr90_48_reg [51]),
        .O(adr_reg_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_42
       (.CI(adr_reg_i_52_n_0),
        .CO({adr_reg_i_42_n_0,adr_reg_i_42_n_1,adr_reg_i_42_n_2,adr_reg_i_42_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr_48_reg [43:42],\<const0>__0__0 ,\<const0>__0__0 }),
        .S({adr_reg_i_53_n_0,adr_reg_i_54_n_0,\I_1/ctr_48_reg [41:40]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_43
       (.I0(\I_1/ctr_48_reg [47]),
        .O(adr_reg_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_44
       (.I0(\I_1/ctr_48_reg [46]),
        .O(adr_reg_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_45
       (.I0(\I_1/ctr_48_reg [45]),
        .O(adr_reg_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_47
       (.CI(adr_reg_i_57_n_0),
        .CO({adr_reg_i_47_n_0,adr_reg_i_47_n_1,adr_reg_i_47_n_2,adr_reg_i_47_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr90_48_reg [43:42],\<const0>__0__0 ,\<const0>__0__0 }),
        .S({adr_reg_i_58_n_0,adr_reg_i_59_n_0,\I_1/ctr90_48_reg [41:40]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_48
       (.I0(\I_1/ctr90_48_reg [47]),
        .O(adr_reg_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_49
       (.I0(\I_1/ctr90_48_reg [46]),
        .O(adr_reg_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_50
       (.I0(\I_1/ctr90_48_reg [45]),
        .O(adr_reg_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_52
       (.CI(adr_reg_i_62_n_0),
        .CO({adr_reg_i_52_n_0,adr_reg_i_52_n_1,adr_reg_i_52_n_2,adr_reg_i_52_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr_48_reg [39:37],\<const0>__0__0 }),
        .S({adr_reg_i_63_n_0,adr_reg_i_64_n_0,adr_reg_i_65_n_0,\I_1/ctr_48_reg [36]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_53
       (.I0(\I_1/ctr_48_reg [43]),
        .O(adr_reg_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_54
       (.I0(\I_1/ctr_48_reg [42]),
        .O(adr_reg_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_57
       (.CI(adr_reg_i_67_n_0),
        .CO({adr_reg_i_57_n_0,adr_reg_i_57_n_1,adr_reg_i_57_n_2,adr_reg_i_57_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\I_1/ctr90_48_reg [39:37],\<const0>__0__0 }),
        .S({adr_reg_i_68_n_0,adr_reg_i_69_n_0,adr_reg_i_70_n_0,\I_1/ctr90_48_reg [36]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_58
       (.I0(\I_1/ctr90_48_reg [43]),
        .O(adr_reg_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_59
       (.I0(\I_1/ctr90_48_reg [42]),
        .O(adr_reg_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_62
       (.CI(adr_reg_i_72_n_0),
        .CO({adr_reg_i_62_n_0,adr_reg_i_62_n_1,adr_reg_i_62_n_2,adr_reg_i_62_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S(\I_1/ctr_48_reg [35:32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_63
       (.I0(\I_1/ctr_48_reg [39]),
        .O(adr_reg_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_64
       (.I0(\I_1/ctr_48_reg [38]),
        .O(adr_reg_i_64_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_65
       (.I0(\I_1/ctr_48_reg [37]),
        .O(adr_reg_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_67
       (.CI(adr_reg_i_77_n_0),
        .CO({adr_reg_i_67_n_0,adr_reg_i_67_n_1,adr_reg_i_67_n_2,adr_reg_i_67_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S(\I_1/ctr90_48_reg [35:32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_68
       (.I0(\I_1/ctr90_48_reg [39]),
        .O(adr_reg_i_68_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_69
       (.I0(\I_1/ctr90_48_reg [38]),
        .O(adr_reg_i_69_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_70
       (.I0(\I_1/ctr90_48_reg [37]),
        .O(adr_reg_i_70_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_72
       (.CI(adr_reg_i_82_n_0),
        .CO({adr_reg_i_72_n_0,adr_reg_i_72_n_1,adr_reg_i_72_n_2,adr_reg_i_72_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr_48_reg [30],\<const0>__0__0 ,\I_1/ctr_48_reg [28]}),
        .S({\I_1/ctr_48_reg [31],adr_reg_i_84_n_0,\I_1/ctr_48_reg [29],adr_reg_i_86_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_77
       (.CI(adr_reg_i_87_n_0),
        .CO({adr_reg_i_77_n_0,adr_reg_i_77_n_1,adr_reg_i_77_n_2,adr_reg_i_77_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\I_1/ctr90_48_reg [30],\<const0>__0__0 ,\I_1/ctr90_48_reg [28]}),
        .S({\I_1/ctr90_48_reg [31],adr_reg_i_89_n_0,\I_1/ctr90_48_reg [29],adr_reg_i_91_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_82
       (.CI(adr_reg_i_92_n_0),
        .CO({adr_reg_i_82_n_0,adr_reg_i_82_n_1,adr_reg_i_82_n_2,adr_reg_i_82_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [25:24]}),
        .S({\I_1/ctr_48_reg [27:26],adr_reg_i_95_n_0,adr_reg_i_96_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_84
       (.I0(\I_1/ctr_48_reg [30]),
        .O(adr_reg_i_84_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_86
       (.I0(\I_1/ctr_48_reg [28]),
        .O(adr_reg_i_86_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_87
       (.CI(adr_reg_i_97_n_0),
        .CO({adr_reg_i_87_n_0,adr_reg_i_87_n_1,adr_reg_i_87_n_2,adr_reg_i_87_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [25:24]}),
        .S({\I_1/ctr90_48_reg [27:26],adr_reg_i_100_n_0,adr_reg_i_101_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_89
       (.I0(\I_1/ctr90_48_reg [30]),
        .O(adr_reg_i_89_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_91
       (.I0(\I_1/ctr90_48_reg [28]),
        .O(adr_reg_i_91_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_92
       (.CI(adr_reg_i_102_n_0),
        .CO({adr_reg_i_92_n_0,adr_reg_i_92_n_1,adr_reg_i_92_n_2,adr_reg_i_92_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr_48_reg [20]}),
        .S({\I_1/ctr_48_reg [23:21],adr_reg_i_106_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_95
       (.I0(\I_1/ctr_48_reg [25]),
        .O(adr_reg_i_95_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    adr_reg_i_96
       (.I0(\I_1/ctr_48_reg [24]),
        .O(adr_reg_i_96_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 adr_reg_i_97
       (.CI(adr_reg_i_107_n_0),
        .CO({adr_reg_i_97_n_0,adr_reg_i_97_n_1,adr_reg_i_97_n_2,adr_reg_i_97_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_1/ctr90_48_reg [20]}),
        .S({\I_1/ctr90_48_reg [23:21],adr_reg_i_111_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hC5)) 
    austastung_i_1
       (.I0(\I_0/i_austastung ),
        .I1(i_austastung_i_3_n_0),
        .I2(\I_0/hlctr0 ),
        .O(austastung_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[13]_i_2 
       (.I0(\I_1/ctr90_48_reg [16]),
        .O(ctr90_48));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[13]_i_4 
       (.I0(\I_1/ctr90_48_reg [14]),
        .O(\ctr90_48[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[13]_i_5 
       (.I0(\I_1/ctr90_48_reg [13]),
        .O(\ctr90_48[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[17]_i_2 
       (.I0(\I_1/ctr90_48_reg [20]),
        .O(\ctr90_48[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[1]_i_2 
       (.I0(\I_1/ctr90_48_reg [4]),
        .O(\ctr90_48[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[1]_i_5 
       (.I0(\I_1/ctr90_48_reg [1]),
        .O(\ctr90_48[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[21]_i_2 
       (.I0(\I_1/ctr90_48_reg [24]),
        .O(\ctr90_48[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[25]_i_2 
       (.I0(\I_1/ctr90_48_reg [28]),
        .O(\ctr90_48[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[25]_i_5 
       (.I0(\I_1/ctr90_48_reg [25]),
        .O(\ctr90_48[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[29]_i_4 
       (.I0(\I_1/ctr90_48_reg [30]),
        .O(\ctr90_48[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[37]_i_3 
       (.I0(\I_1/ctr90_48_reg [39]),
        .O(\ctr90_48[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[37]_i_4 
       (.I0(\I_1/ctr90_48_reg [38]),
        .O(\ctr90_48[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[37]_i_5 
       (.I0(\I_1/ctr90_48_reg [37]),
        .O(\ctr90_48[37]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[41]_i_3 
       (.I0(\I_1/ctr90_48_reg [43]),
        .O(\ctr90_48[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[41]_i_4 
       (.I0(\I_1/ctr90_48_reg [42]),
        .O(\ctr90_48[41]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[45]_i_3 
       (.I0(\I_1/ctr90_48_reg [47]),
        .O(\ctr90_48[45]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[45]_i_4 
       (.I0(\I_1/ctr90_48_reg [46]),
        .O(\ctr90_48[45]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[45]_i_5 
       (.I0(\I_1/ctr90_48_reg [45]),
        .O(\ctr90_48[45]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[49]_i_2 
       (.I0(\I_1/ctr90_48_reg [52]),
        .O(\ctr90_48[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[49]_i_3 
       (.I0(\I_1/ctr90_48_reg [51]),
        .O(\ctr90_48[49]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[53]_i_2 
       (.I0(\I_1/ctr90_48_reg [56]),
        .O(\ctr90_48[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[53]_i_5 
       (.I0(\I_1/ctr90_48_reg [53]),
        .O(\ctr90_48[53]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[57]_i_2 
       (.I0(\I_1/ctr90_48_reg [60]),
        .O(\ctr90_48[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[57]_i_3 
       (.I0(\I_1/ctr90_48_reg [59]),
        .O(\ctr90_48[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[5]_i_3 
       (.I0(\I_1/ctr90_48_reg [7]),
        .O(\ctr90_48[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[5]_i_4 
       (.I0(\I_1/ctr90_48_reg [6]),
        .O(\ctr90_48[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[5]_i_5 
       (.I0(\I_1/ctr90_48_reg [5]),
        .O(\ctr90_48[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[9]_i_2 
       (.I0(\I_1/ctr90_48_reg [12]),
        .O(\ctr90_48[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr90_48[9]_i_4 
       (.I0(\I_1/ctr90_48_reg [10]),
        .O(\ctr90_48[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[13]_i_1 
       (.CI(\ctr90_48_reg[9]_i_1_n_0 ),
        .CO(ctr90_48_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[13]_i_1_n_4 ,\ctr90_48_reg[13]_i_1_n_5 ,\ctr90_48_reg[13]_i_1_n_6 ,\ctr90_48_reg[13]_i_1_n_7 }),
        .S({ctr90_48,\I_1/ctr90_48_reg [15],\ctr90_48[13]_i_4_n_0 ,\ctr90_48[13]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[17]_i_1 
       (.CI(ctr90_48_reg[3]),
        .CO({\ctr90_48_reg[17]_i_1_n_0 ,\ctr90_48_reg[17]_i_1_n_1 ,\ctr90_48_reg[17]_i_1_n_2 ,\ctr90_48_reg[17]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[17]_i_1_n_4 ,\ctr90_48_reg[17]_i_1_n_5 ,\ctr90_48_reg[17]_i_1_n_6 ,\ctr90_48_reg[17]_i_1_n_7 }),
        .S({\ctr90_48[17]_i_2_n_0 ,\I_1/ctr90_48_reg [19:17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[1]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\ctr90_48_reg[1]_i_1_n_0 ,\ctr90_48_reg[1]_i_1_n_1 ,\ctr90_48_reg[1]_i_1_n_2 ,\ctr90_48_reg[1]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[1]_i_1_n_4 ,\ctr90_48_reg[1]_i_1_n_5 ,\ctr90_48_reg[1]_i_1_n_6 ,\ctr90_48_reg[1]_i_1_n_7 }),
        .S({\ctr90_48[1]_i_2_n_0 ,\I_1/ctr90_48_reg [3:2],\ctr90_48[1]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[21]_i_1 
       (.CI(\ctr90_48_reg[17]_i_1_n_0 ),
        .CO({\ctr90_48_reg[21]_i_1_n_0 ,\ctr90_48_reg[21]_i_1_n_1 ,\ctr90_48_reg[21]_i_1_n_2 ,\ctr90_48_reg[21]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[21]_i_1_n_4 ,\ctr90_48_reg[21]_i_1_n_5 ,\ctr90_48_reg[21]_i_1_n_6 ,\ctr90_48_reg[21]_i_1_n_7 }),
        .S({\ctr90_48[21]_i_2_n_0 ,\I_1/ctr90_48_reg [23:21]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[25]_i_1 
       (.CI(\ctr90_48_reg[21]_i_1_n_0 ),
        .CO({\ctr90_48_reg[25]_i_1_n_0 ,\ctr90_48_reg[25]_i_1_n_1 ,\ctr90_48_reg[25]_i_1_n_2 ,\ctr90_48_reg[25]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[25]_i_1_n_4 ,\ctr90_48_reg[25]_i_1_n_5 ,\ctr90_48_reg[25]_i_1_n_6 ,\ctr90_48_reg[25]_i_1_n_7 }),
        .S({\ctr90_48[25]_i_2_n_0 ,\I_1/ctr90_48_reg [27:26],\ctr90_48[25]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[29]_i_1 
       (.CI(\ctr90_48_reg[25]_i_1_n_0 ),
        .CO({\ctr90_48_reg[29]_i_1_n_0 ,\ctr90_48_reg[29]_i_1_n_1 ,\ctr90_48_reg[29]_i_1_n_2 ,\ctr90_48_reg[29]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[29]_i_1_n_4 ,\ctr90_48_reg[29]_i_1_n_5 ,\ctr90_48_reg[29]_i_1_n_6 ,\ctr90_48_reg[29]_i_1_n_7 }),
        .S({\I_1/ctr90_48_reg [32:31],\ctr90_48[29]_i_4_n_0 ,\I_1/ctr90_48_reg [29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[33]_i_1 
       (.CI(\ctr90_48_reg[29]_i_1_n_0 ),
        .CO({\ctr90_48_reg[33]_i_1_n_0 ,\ctr90_48_reg[33]_i_1_n_1 ,\ctr90_48_reg[33]_i_1_n_2 ,\ctr90_48_reg[33]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[33]_i_1_n_4 ,\ctr90_48_reg[33]_i_1_n_5 ,\ctr90_48_reg[33]_i_1_n_6 ,\ctr90_48_reg[33]_i_1_n_7 }),
        .S(\I_1/ctr90_48_reg [36:33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[37]_i_1 
       (.CI(\ctr90_48_reg[33]_i_1_n_0 ),
        .CO({\ctr90_48_reg[37]_i_1_n_0 ,\ctr90_48_reg[37]_i_1_n_1 ,\ctr90_48_reg[37]_i_1_n_2 ,\ctr90_48_reg[37]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[37]_i_1_n_4 ,\ctr90_48_reg[37]_i_1_n_5 ,\ctr90_48_reg[37]_i_1_n_6 ,\ctr90_48_reg[37]_i_1_n_7 }),
        .S({\I_1/ctr90_48_reg [40],\ctr90_48[37]_i_3_n_0 ,\ctr90_48[37]_i_4_n_0 ,\ctr90_48[37]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[41]_i_1 
       (.CI(\ctr90_48_reg[37]_i_1_n_0 ),
        .CO({\ctr90_48_reg[41]_i_1_n_0 ,\ctr90_48_reg[41]_i_1_n_1 ,\ctr90_48_reg[41]_i_1_n_2 ,\ctr90_48_reg[41]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[41]_i_1_n_4 ,\ctr90_48_reg[41]_i_1_n_5 ,\ctr90_48_reg[41]_i_1_n_6 ,\ctr90_48_reg[41]_i_1_n_7 }),
        .S({\I_1/ctr90_48_reg [44],\ctr90_48[41]_i_3_n_0 ,\ctr90_48[41]_i_4_n_0 ,\I_1/ctr90_48_reg [41]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[45]_i_1 
       (.CI(\ctr90_48_reg[41]_i_1_n_0 ),
        .CO({\ctr90_48_reg[45]_i_1_n_0 ,\ctr90_48_reg[45]_i_1_n_1 ,\ctr90_48_reg[45]_i_1_n_2 ,\ctr90_48_reg[45]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[45]_i_1_n_4 ,\ctr90_48_reg[45]_i_1_n_5 ,\ctr90_48_reg[45]_i_1_n_6 ,\ctr90_48_reg[45]_i_1_n_7 }),
        .S({\I_1/ctr90_48_reg [48],\ctr90_48[45]_i_3_n_0 ,\ctr90_48[45]_i_4_n_0 ,\ctr90_48[45]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[49]_i_1 
       (.CI(\ctr90_48_reg[45]_i_1_n_0 ),
        .CO({\ctr90_48_reg[49]_i_1_n_0 ,\ctr90_48_reg[49]_i_1_n_1 ,\ctr90_48_reg[49]_i_1_n_2 ,\ctr90_48_reg[49]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[49]_i_1_n_4 ,\ctr90_48_reg[49]_i_1_n_5 ,\ctr90_48_reg[49]_i_1_n_6 ,\ctr90_48_reg[49]_i_1_n_7 }),
        .S({\ctr90_48[49]_i_2_n_0 ,\ctr90_48[49]_i_3_n_0 ,\I_1/ctr90_48_reg [50:49]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[53]_i_1 
       (.CI(\ctr90_48_reg[49]_i_1_n_0 ),
        .CO({\ctr90_48_reg[53]_i_1_n_0 ,\ctr90_48_reg[53]_i_1_n_1 ,\ctr90_48_reg[53]_i_1_n_2 ,\ctr90_48_reg[53]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[53]_i_1_n_4 ,\ctr90_48_reg[53]_i_1_n_5 ,\ctr90_48_reg[53]_i_1_n_6 ,\ctr90_48_reg[53]_i_1_n_7 }),
        .S({\ctr90_48[53]_i_2_n_0 ,\I_1/ctr90_48_reg [55:54],\ctr90_48[53]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[57]_i_1 
       (.CI(\ctr90_48_reg[53]_i_1_n_0 ),
        .CO({\ctr90_48_reg[57]_i_1_n_0 ,\ctr90_48_reg[57]_i_1_n_1 ,\ctr90_48_reg[57]_i_1_n_2 ,\ctr90_48_reg[57]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[57]_i_1_n_4 ,\ctr90_48_reg[57]_i_1_n_5 ,\ctr90_48_reg[57]_i_1_n_6 ,\ctr90_48_reg[57]_i_1_n_7 }),
        .S({\ctr90_48[57]_i_2_n_0 ,\ctr90_48[57]_i_3_n_0 ,\I_1/ctr90_48_reg [58:57]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[5]_i_1 
       (.CI(\ctr90_48_reg[1]_i_1_n_0 ),
        .CO({\ctr90_48_reg[5]_i_1_n_0 ,\ctr90_48_reg[5]_i_1_n_1 ,\ctr90_48_reg[5]_i_1_n_2 ,\ctr90_48_reg[5]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr90_48_reg[5]_i_1_n_4 ,\ctr90_48_reg[5]_i_1_n_5 ,\ctr90_48_reg[5]_i_1_n_6 ,\ctr90_48_reg[5]_i_1_n_7 }),
        .S({\I_1/ctr90_48_reg [8],\ctr90_48[5]_i_3_n_0 ,\ctr90_48[5]_i_4_n_0 ,\ctr90_48[5]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[61]_i_1 
       (.CI(\ctr90_48_reg[57]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[61]_i_1_n_4 ,\ctr90_48_reg[61]_i_1_n_5 ,\ctr90_48_reg[61]_i_1_n_6 ,\ctr90_48_reg[61]_i_1_n_7 }),
        .S({\<const0>__0__0 ,\I_1/ctr90_48_reg [63:61]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr90_48_reg[9]_i_1 
       (.CI(\ctr90_48_reg[5]_i_1_n_0 ),
        .CO({\ctr90_48_reg[9]_i_1_n_0 ,\ctr90_48_reg[9]_i_1_n_1 ,\ctr90_48_reg[9]_i_1_n_2 ,\ctr90_48_reg[9]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr90_48_reg[9]_i_1_n_4 ,\ctr90_48_reg[9]_i_1_n_5 ,\ctr90_48_reg[9]_i_1_n_6 ,\ctr90_48_reg[9]_i_1_n_7 }),
        .S({\ctr90_48[9]_i_2_n_0 ,\I_1/ctr90_48_reg [11],\ctr90_48[9]_i_4_n_0 ,\I_1/ctr90_48_reg [9]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[13]_i_2 
       (.I0(\I_1/ctr_48_reg [16]),
        .O(ctr_48));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[13]_i_4 
       (.I0(\I_1/ctr_48_reg [14]),
        .O(\ctr_48[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[13]_i_5 
       (.I0(\I_1/ctr_48_reg [13]),
        .O(\ctr_48[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[17]_i_2 
       (.I0(\I_1/ctr_48_reg [20]),
        .O(\ctr_48[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[1]_i_2 
       (.I0(\I_1/ctr_48_reg [4]),
        .O(\ctr_48[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[1]_i_5 
       (.I0(\I_1/ctr_48_reg [1]),
        .O(\ctr_48[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[21]_i_2 
       (.I0(\I_1/ctr_48_reg [24]),
        .O(\ctr_48[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[25]_i_2 
       (.I0(\I_1/ctr_48_reg [28]),
        .O(\ctr_48[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[25]_i_5 
       (.I0(\I_1/ctr_48_reg [25]),
        .O(\ctr_48[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[29]_i_4 
       (.I0(\I_1/ctr_48_reg [30]),
        .O(\ctr_48[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[37]_i_3 
       (.I0(\I_1/ctr_48_reg [39]),
        .O(\ctr_48[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[37]_i_4 
       (.I0(\I_1/ctr_48_reg [38]),
        .O(\ctr_48[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[37]_i_5 
       (.I0(\I_1/ctr_48_reg [37]),
        .O(\ctr_48[37]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[41]_i_3 
       (.I0(\I_1/ctr_48_reg [43]),
        .O(\ctr_48[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[41]_i_4 
       (.I0(\I_1/ctr_48_reg [42]),
        .O(\ctr_48[41]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[45]_i_3 
       (.I0(\I_1/ctr_48_reg [47]),
        .O(\ctr_48[45]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[45]_i_4 
       (.I0(\I_1/ctr_48_reg [46]),
        .O(\ctr_48[45]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[45]_i_5 
       (.I0(\I_1/ctr_48_reg [45]),
        .O(\ctr_48[45]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[49]_i_2 
       (.I0(\I_1/ctr_48_reg [52]),
        .O(\ctr_48[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[49]_i_3 
       (.I0(\I_1/ctr_48_reg [51]),
        .O(\ctr_48[49]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[53]_i_2 
       (.I0(\I_1/ctr_48_reg [56]),
        .O(\ctr_48[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[53]_i_5 
       (.I0(\I_1/ctr_48_reg [53]),
        .O(\ctr_48[53]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[57]_i_2 
       (.I0(\I_1/ctr_48_reg [60]),
        .O(\ctr_48[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[57]_i_3 
       (.I0(\I_1/ctr_48_reg [59]),
        .O(\ctr_48[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[5]_i_3 
       (.I0(\I_1/ctr_48_reg [7]),
        .O(\ctr_48[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[5]_i_4 
       (.I0(\I_1/ctr_48_reg [6]),
        .O(\ctr_48[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[5]_i_5 
       (.I0(\I_1/ctr_48_reg [5]),
        .O(\ctr_48[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[9]_i_2 
       (.I0(\I_1/ctr_48_reg [12]),
        .O(\ctr_48[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \ctr_48[9]_i_4 
       (.I0(\I_1/ctr_48_reg [10]),
        .O(\ctr_48[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[13]_i_1 
       (.CI(\ctr_48_reg[9]_i_1_n_0 ),
        .CO(ctr_48_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[13]_i_1_n_4 ,\ctr_48_reg[13]_i_1_n_5 ,\ctr_48_reg[13]_i_1_n_6 ,\ctr_48_reg[13]_i_1_n_7 }),
        .S({ctr_48,\I_1/ctr_48_reg [15],\ctr_48[13]_i_4_n_0 ,\ctr_48[13]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[17]_i_1 
       (.CI(ctr_48_reg[3]),
        .CO({\ctr_48_reg[17]_i_1_n_0 ,\ctr_48_reg[17]_i_1_n_1 ,\ctr_48_reg[17]_i_1_n_2 ,\ctr_48_reg[17]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[17]_i_1_n_4 ,\ctr_48_reg[17]_i_1_n_5 ,\ctr_48_reg[17]_i_1_n_6 ,\ctr_48_reg[17]_i_1_n_7 }),
        .S({\ctr_48[17]_i_2_n_0 ,\I_1/ctr_48_reg [19:17]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[1]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\ctr_48_reg[1]_i_1_n_0 ,\ctr_48_reg[1]_i_1_n_1 ,\ctr_48_reg[1]_i_1_n_2 ,\ctr_48_reg[1]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[1]_i_1_n_4 ,\ctr_48_reg[1]_i_1_n_5 ,\ctr_48_reg[1]_i_1_n_6 ,\ctr_48_reg[1]_i_1_n_7 }),
        .S({\ctr_48[1]_i_2_n_0 ,\I_1/ctr_48_reg [3:2],\ctr_48[1]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[21]_i_1 
       (.CI(\ctr_48_reg[17]_i_1_n_0 ),
        .CO({\ctr_48_reg[21]_i_1_n_0 ,\ctr_48_reg[21]_i_1_n_1 ,\ctr_48_reg[21]_i_1_n_2 ,\ctr_48_reg[21]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[21]_i_1_n_4 ,\ctr_48_reg[21]_i_1_n_5 ,\ctr_48_reg[21]_i_1_n_6 ,\ctr_48_reg[21]_i_1_n_7 }),
        .S({\ctr_48[21]_i_2_n_0 ,\I_1/ctr_48_reg [23:21]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[25]_i_1 
       (.CI(\ctr_48_reg[21]_i_1_n_0 ),
        .CO({\ctr_48_reg[25]_i_1_n_0 ,\ctr_48_reg[25]_i_1_n_1 ,\ctr_48_reg[25]_i_1_n_2 ,\ctr_48_reg[25]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[25]_i_1_n_4 ,\ctr_48_reg[25]_i_1_n_5 ,\ctr_48_reg[25]_i_1_n_6 ,\ctr_48_reg[25]_i_1_n_7 }),
        .S({\ctr_48[25]_i_2_n_0 ,\I_1/ctr_48_reg [27:26],\ctr_48[25]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[29]_i_1 
       (.CI(\ctr_48_reg[25]_i_1_n_0 ),
        .CO({\ctr_48_reg[29]_i_1_n_0 ,\ctr_48_reg[29]_i_1_n_1 ,\ctr_48_reg[29]_i_1_n_2 ,\ctr_48_reg[29]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[29]_i_1_n_4 ,\ctr_48_reg[29]_i_1_n_5 ,\ctr_48_reg[29]_i_1_n_6 ,\ctr_48_reg[29]_i_1_n_7 }),
        .S({\I_1/ctr_48_reg [32:31],\ctr_48[29]_i_4_n_0 ,\I_1/ctr_48_reg [29]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[33]_i_1 
       (.CI(\ctr_48_reg[29]_i_1_n_0 ),
        .CO({\ctr_48_reg[33]_i_1_n_0 ,\ctr_48_reg[33]_i_1_n_1 ,\ctr_48_reg[33]_i_1_n_2 ,\ctr_48_reg[33]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[33]_i_1_n_4 ,\ctr_48_reg[33]_i_1_n_5 ,\ctr_48_reg[33]_i_1_n_6 ,\ctr_48_reg[33]_i_1_n_7 }),
        .S(\I_1/ctr_48_reg [36:33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[37]_i_1 
       (.CI(\ctr_48_reg[33]_i_1_n_0 ),
        .CO({\ctr_48_reg[37]_i_1_n_0 ,\ctr_48_reg[37]_i_1_n_1 ,\ctr_48_reg[37]_i_1_n_2 ,\ctr_48_reg[37]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[37]_i_1_n_4 ,\ctr_48_reg[37]_i_1_n_5 ,\ctr_48_reg[37]_i_1_n_6 ,\ctr_48_reg[37]_i_1_n_7 }),
        .S({\I_1/ctr_48_reg [40],\ctr_48[37]_i_3_n_0 ,\ctr_48[37]_i_4_n_0 ,\ctr_48[37]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[41]_i_1 
       (.CI(\ctr_48_reg[37]_i_1_n_0 ),
        .CO({\ctr_48_reg[41]_i_1_n_0 ,\ctr_48_reg[41]_i_1_n_1 ,\ctr_48_reg[41]_i_1_n_2 ,\ctr_48_reg[41]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[41]_i_1_n_4 ,\ctr_48_reg[41]_i_1_n_5 ,\ctr_48_reg[41]_i_1_n_6 ,\ctr_48_reg[41]_i_1_n_7 }),
        .S({\I_1/ctr_48_reg [44],\ctr_48[41]_i_3_n_0 ,\ctr_48[41]_i_4_n_0 ,\I_1/ctr_48_reg [41]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[45]_i_1 
       (.CI(\ctr_48_reg[41]_i_1_n_0 ),
        .CO({\ctr_48_reg[45]_i_1_n_0 ,\ctr_48_reg[45]_i_1_n_1 ,\ctr_48_reg[45]_i_1_n_2 ,\ctr_48_reg[45]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[45]_i_1_n_4 ,\ctr_48_reg[45]_i_1_n_5 ,\ctr_48_reg[45]_i_1_n_6 ,\ctr_48_reg[45]_i_1_n_7 }),
        .S({\I_1/ctr_48_reg [48],\ctr_48[45]_i_3_n_0 ,\ctr_48[45]_i_4_n_0 ,\ctr_48[45]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[49]_i_1 
       (.CI(\ctr_48_reg[45]_i_1_n_0 ),
        .CO({\ctr_48_reg[49]_i_1_n_0 ,\ctr_48_reg[49]_i_1_n_1 ,\ctr_48_reg[49]_i_1_n_2 ,\ctr_48_reg[49]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[49]_i_1_n_4 ,\ctr_48_reg[49]_i_1_n_5 ,\ctr_48_reg[49]_i_1_n_6 ,\ctr_48_reg[49]_i_1_n_7 }),
        .S({\ctr_48[49]_i_2_n_0 ,\ctr_48[49]_i_3_n_0 ,\I_1/ctr_48_reg [50:49]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[53]_i_1 
       (.CI(\ctr_48_reg[49]_i_1_n_0 ),
        .CO({\ctr_48_reg[53]_i_1_n_0 ,\ctr_48_reg[53]_i_1_n_1 ,\ctr_48_reg[53]_i_1_n_2 ,\ctr_48_reg[53]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[53]_i_1_n_4 ,\ctr_48_reg[53]_i_1_n_5 ,\ctr_48_reg[53]_i_1_n_6 ,\ctr_48_reg[53]_i_1_n_7 }),
        .S({\ctr_48[53]_i_2_n_0 ,\I_1/ctr_48_reg [55:54],\ctr_48[53]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[57]_i_1 
       (.CI(\ctr_48_reg[53]_i_1_n_0 ),
        .CO({\ctr_48_reg[57]_i_1_n_0 ,\ctr_48_reg[57]_i_1_n_1 ,\ctr_48_reg[57]_i_1_n_2 ,\ctr_48_reg[57]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[57]_i_1_n_4 ,\ctr_48_reg[57]_i_1_n_5 ,\ctr_48_reg[57]_i_1_n_6 ,\ctr_48_reg[57]_i_1_n_7 }),
        .S({\ctr_48[57]_i_2_n_0 ,\ctr_48[57]_i_3_n_0 ,\I_1/ctr_48_reg [58:57]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[5]_i_1 
       (.CI(\ctr_48_reg[1]_i_1_n_0 ),
        .CO({\ctr_48_reg[5]_i_1_n_0 ,\ctr_48_reg[5]_i_1_n_1 ,\ctr_48_reg[5]_i_1_n_2 ,\ctr_48_reg[5]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\ctr_48_reg[5]_i_1_n_4 ,\ctr_48_reg[5]_i_1_n_5 ,\ctr_48_reg[5]_i_1_n_6 ,\ctr_48_reg[5]_i_1_n_7 }),
        .S({\I_1/ctr_48_reg [8],\ctr_48[5]_i_3_n_0 ,\ctr_48[5]_i_4_n_0 ,\ctr_48[5]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[61]_i_1 
       (.CI(\ctr_48_reg[57]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[61]_i_1_n_4 ,\ctr_48_reg[61]_i_1_n_5 ,\ctr_48_reg[61]_i_1_n_6 ,\ctr_48_reg[61]_i_1_n_7 }),
        .S({\<const0>__0__0 ,\I_1/ctr_48_reg [63:61]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \ctr_48_reg[9]_i_1 
       (.CI(\ctr_48_reg[5]_i_1_n_0 ),
        .CO({\ctr_48_reg[9]_i_1_n_0 ,\ctr_48_reg[9]_i_1_n_1 ,\ctr_48_reg[9]_i_1_n_2 ,\ctr_48_reg[9]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 }),
        .O({\ctr_48_reg[9]_i_1_n_4 ,\ctr_48_reg[9]_i_1_n_5 ,\ctr_48_reg[9]_i_1_n_6 ,\ctr_48_reg[9]_i_1_n_7 }),
        .S({\ctr_48[9]_i_2_n_0 ,\I_1/ctr_48_reg [11],\ctr_48[9]_i_4_n_0 ,\I_1/ctr_48_reg [9]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[12]_i_2 
       (.CI(\data_reg[8]_i_2_n_0 ),
        .CO({\data_reg[12]_i_2_n_0 ,\data_reg[12]_i_2_n_1 ,\data_reg[12]_i_2_n_2 ,\data_reg[12]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(data0[12:9]),
        .S({\I_2/data ,\I_2/data[12]_i_4_n_0 ,\I_2/data[12]_i_5_n_0 ,\I_2/data[12]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[12]_i_2__0 
       (.CI(\data_reg[8]_i_2__0_n_0 ),
        .CO(data_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\data_reg[12]_i_2__0_n_4 ,\data_reg[12]_i_2__0_n_5 ,\data_reg[12]_i_2__0_n_6 ,\data_reg[12]_i_2__0_n_7 }),
        .S({\I_1/data[12]_i_3_n_0 ,\I_1/data[12]_i_4_n_0 ,\I_1/data[12]_i_5_n_0 ,\I_1/data[12]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[15]_i_2 
       (.CI(\data_reg[12]_i_2_n_0 ),
        .CO({\data_reg[15]_i_2_n_0 ,\data_reg[15]_i_2_n_1 ,\data_reg[15]_i_2_n_2 ,\data_reg[15]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\data_reg[15]_i_2_n_4 ,\data_reg[15]_i_2_n_5 ,data0[14:13]}),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\I_2/data[15]_i_3_n_0 ,\I_2/data[15]_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[15]_i_2__0 
       (.CI(data_reg[3]),
        .CO({\data_reg[15]_i_2__0_n_0 ,\data_reg[15]_i_2__0_n_1 ,\data_reg[15]_i_2__0_n_2 ,\data_reg[15]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\data_reg[15]_i_2__0_n_4 ,\data_reg[15]_i_2__0_n_5 ,\data_reg[15]_i_2__0_n_6 ,\data_reg[15]_i_2__0_n_7 }),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\I_1/data[15]_i_3_n_0 ,\I_1/data[15]_i_4_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[4]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\data_reg[4]_i_2_n_0 ,\data_reg[4]_i_2_n_1 ,\data_reg[4]_i_2_n_2 ,\data_reg[4]_i_2_n_3 }),
        .CYINIT(\I_2/data[4]_i_3_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(data0[4:1]),
        .S({\I_2/data[4]_i_4_n_0 ,\I_2/data[4]_i_5_n_0 ,\I_2/data[4]_i_6_n_0 ,\I_2/data[4]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[4]_i_2__0 
       (.CI(\<const0>__0__0 ),
        .CO({\data_reg[4]_i_2__0_n_0 ,\data_reg[4]_i_2__0_n_1 ,\data_reg[4]_i_2__0_n_2 ,\data_reg[4]_i_2__0_n_3 }),
        .CYINIT(\I_1/data[4]_i_3_n_0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\data_reg[4]_i_2__0_n_4 ,\data_reg[4]_i_2__0_n_5 ,\data_reg[4]_i_2__0_n_6 ,\data_reg[4]_i_2__0_n_7 }),
        .S({\I_1/data[4]_i_4_n_0 ,\I_1/data[4]_i_5_n_0 ,\I_1/data[4]_i_6_n_0 ,\I_1/data[4]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[8]_i_2 
       (.CI(\data_reg[4]_i_2_n_0 ),
        .CO({\data_reg[8]_i_2_n_0 ,\data_reg[8]_i_2_n_1 ,\data_reg[8]_i_2_n_2 ,\data_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(data0[8:5]),
        .S({\I_2/data[8]_i_3_n_0 ,\I_2/data[8]_i_4_n_0 ,\I_2/data[8]_i_5_n_0 ,\I_2/data[8]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \data_reg[8]_i_2__0 
       (.CI(\data_reg[4]_i_2__0_n_0 ),
        .CO({\data_reg[8]_i_2__0_n_0 ,\data_reg[8]_i_2__0_n_1 ,\data_reg[8]_i_2__0_n_2 ,\data_reg[8]_i_2__0_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\data_reg[8]_i_2__0_n_4 ,\data_reg[8]_i_2__0_n_5 ,\data_reg[8]_i_2__0_n_6 ,\data_reg[8]_i_2__0_n_7 }),
        .S({\I_1/data[8]_i_3_n_0 ,\I_1/data[8]_i_4_n_0 ,\I_1/data[8]_i_5_n_0 ,\I_1/data[8]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__0_i_1
       (.I0(\I_0/pixctr2_carry__2_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_5 ),
        .O(en_bild1_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__0_i_2
       (.I0(\I_0/pixctr2_carry__1_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_7 ),
        .O(en_bild1_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__0_i_3
       (.I0(\I_0/pixctr2_carry__1_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_5 ),
        .O(en_bild1_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__0_i_4
       (.I0(\I_0/pixctr2_carry__0_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(en_bild1_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__0_i_5
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(en_bild1_inferred__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__0_i_6
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(en_bild1_inferred__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__0_i_7
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(en_bild1_inferred__0_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__0_i_8
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(en_bild1_inferred__0_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__1_i_1
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_5 ),
        .O(en_bild1_inferred__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__1_i_2
       (.I0(\I_0/pixctr2_carry__3_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_7 ),
        .O(en_bild1_inferred__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__1_i_3
       (.I0(\I_0/pixctr2_carry__3_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_5 ),
        .O(en_bild1_inferred__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__1_i_4
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_7 ),
        .O(en_bild1_inferred__0_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__1_i_5
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(en_bild1_inferred__0_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__1_i_6
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(en_bild1_inferred__0_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__1_i_7
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(en_bild1_inferred__0_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__1_i_8
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(en_bild1_inferred__0_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild1_inferred__0_carry__2_i_1
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_bild1_inferred__0_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__2_i_2
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__6_n_7 ),
        .O(en_bild1_inferred__0_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__2_i_3
       (.I0(\I_0/pixctr2_carry__5_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_5 ),
        .O(en_bild1_inferred__0_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_bild1_inferred__0_carry__2_i_4
       (.I0(\I_0/pixctr2_carry__4_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_7 ),
        .O(en_bild1_inferred__0_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    en_bild1_inferred__0_carry__2_i_5
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_bild1_inferred__0_carry__2_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__2_i_6
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(en_bild1_inferred__0_carry__2_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__2_i_7
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(en_bild1_inferred__0_carry__2_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild1_inferred__0_carry__2_i_8
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(en_bild1_inferred__0_carry__2_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    en_bild1_inferred__0_carry_i_1
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(en_bild1_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_bild1_inferred__0_carry_i_2
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_bild1_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild1_inferred__0_carry_i_3
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_7 ),
        .I2(\I_0/pixctr_reg_n_0_ ),
        .O(en_bild1_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild1_inferred__0_carry_i_4
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(en_bild1_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    en_bild1_inferred__0_carry_i_5
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(en_bild1_inferred__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    en_bild1_inferred__0_carry_i_6
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(en_bild1_inferred__0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    en_bild1_inferred__0_carry_i_7
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(en_bild1_inferred__0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    en_bild_i_1
       (.I0(\I_0/en_bild1 ),
        .I1(\I_0/en_bild12_in ),
        .O(\I_0/en_bild0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_11
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(en_bild_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_12
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(en_bild_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_13
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(en_bild_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_14
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(en_bild_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    en_bild_i_16
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_bild_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_17
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(en_bild_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_18
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(en_bild_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_19
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(en_bild_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    en_bild_i_2
       (.I0(reset),
        .O(en_bild_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    en_bild_i_20
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(en_bild_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    en_bild_i_21
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .O(en_bild_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    en_bild_i_22
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .O(en_bild_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    en_bild_i_23
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .O(en_bild_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCE)) 
    en_bild_i_24
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(en_bild_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild_i_25
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(en_bild_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild_i_26
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(en_bild_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_bild_i_27
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(en_bild_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    en_bild_i_28
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr_reg_n_0_ ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(en_bild_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_bild_i_5
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_bild_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    en_bild_i_6
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_bild_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_7
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(en_bild_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_8
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(en_bild_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_bild_i_9
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(en_bild_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_bild_reg_i_10
       (.CI(en_bild_reg_i_15_n_0),
        .CO({en_bild_reg_i_10_n_0,en_bild_reg_i_10_n_1,en_bild_reg_i_10_n_2,en_bild_reg_i_10_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,en_bild_i_16_n_0}),
        .S({en_bild_i_17_n_0,en_bild_i_18_n_0,en_bild_i_19_n_0,en_bild_i_20_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_bild_reg_i_15
       (.CI(\<const0>__0__0 ),
        .CO({en_bild_reg_i_15_n_0,en_bild_reg_i_15_n_1,en_bild_reg_i_15_n_2,en_bild_reg_i_15_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({en_bild_i_21_n_0,en_bild_i_22_n_0,en_bild_i_23_n_0,en_bild_i_24_n_0}),
        .S({en_bild_i_25_n_0,en_bild_i_26_n_0,en_bild_i_27_n_0,en_bild_i_28_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_bild_reg_i_3
       (.CI(en_bild_reg_i_4_n_0),
        .CO({\I_0/en_bild1 ,en_bild_reg_i_3_n_1,en_bild_reg_i_3_n_2,en_bild_reg_i_3_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_bild_i_5_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({en_bild_i_6_n_0,en_bild_i_7_n_0,en_bild_i_8_n_0,en_bild_i_9_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_bild_reg_i_4
       (.CI(en_bild_reg_i_10_n_0),
        .CO({en_bild_reg_i_4_n_0,en_bild_reg_i_4_n_1,en_bild_reg_i_4_n_2,en_bild_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({en_bild_i_11_n_0,en_bild_i_12_n_0,en_bild_i_13_n_0,en_bild_i_14_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    en_burst_i_1
       (.I0(\I_0/en_burst1 ),
        .I1(\I_0/en_burst10_in ),
        .O(\I_0/en_burst0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_burst_i_11
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_burst_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_12
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__6_n_7 ),
        .O(en_burst_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_13
       (.I0(\I_0/pixctr2_carry__5_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_5 ),
        .O(en_burst_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_14
       (.I0(\I_0/pixctr2_carry__4_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_7 ),
        .O(en_burst_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    en_burst_i_15
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_burst_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_16
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(en_burst_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_17
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(en_burst_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_18
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(en_burst_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_20
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(en_burst_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_21
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(en_burst_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_22
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(en_burst_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_23
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(en_burst_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_25
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_5 ),
        .O(en_burst_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_26
       (.I0(\I_0/pixctr2_carry__3_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_7 ),
        .O(en_burst_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_27
       (.I0(\I_0/pixctr2_carry__3_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_5 ),
        .O(en_burst_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_28
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_7 ),
        .O(en_burst_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_29
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(en_burst_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_30
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(en_burst_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_31
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(en_burst_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_32
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(en_burst_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_34
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(en_burst_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_35
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(en_burst_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_36
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(en_burst_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_37
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(en_burst_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_39
       (.I0(\I_0/pixctr2_carry__2_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_5 ),
        .O(en_burst_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_40
       (.I0(\I_0/pixctr2_carry__1_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_7 ),
        .O(en_burst_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_41
       (.I0(\I_0/pixctr2_carry__1_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_5 ),
        .O(en_burst_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_42
       (.I0(\I_0/pixctr2_carry__0_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(en_burst_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_43
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(en_burst_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_44
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(en_burst_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_45
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(en_burst_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_46
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(en_burst_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_47
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(en_burst_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    en_burst_i_48
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(en_burst_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_49
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(en_burst_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_burst_i_5
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_burst_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    en_burst_i_50
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_7 ),
        .O(en_burst_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    en_burst_i_51
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(en_burst_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    en_burst_i_52
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(en_burst_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    en_burst_i_53
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_6 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(en_burst_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    en_burst_i_54
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(en_burst_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_burst_i_55
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_burst_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_burst_i_56
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_burst_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    en_burst_i_57
       (.I0(\I_0/pixctr2_carry_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(en_burst_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    en_burst_i_58
       (.I0(\I_0/pixctr2_carry_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(en_burst_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    en_burst_i_59
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(en_burst_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    en_burst_i_6
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(en_burst_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    en_burst_i_60
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(en_burst_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_61
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(en_burst_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    en_burst_i_62
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr_reg_n_0_ ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(en_burst_i_62_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_7
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(en_burst_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_8
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(en_burst_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    en_burst_i_9
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(en_burst_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_10
       (.CI(en_burst_reg_i_24_n_0),
        .CO({en_burst_reg_i_10_n_0,en_burst_reg_i_10_n_1,en_burst_reg_i_10_n_2,en_burst_reg_i_10_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_burst_i_25_n_0,en_burst_i_26_n_0,en_burst_i_27_n_0,en_burst_i_28_n_0}),
        .S({en_burst_i_29_n_0,en_burst_i_30_n_0,en_burst_i_31_n_0,en_burst_i_32_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_19
       (.CI(en_burst_reg_i_33_n_0),
        .CO({en_burst_reg_i_19_n_0,en_burst_reg_i_19_n_1,en_burst_reg_i_19_n_2,en_burst_reg_i_19_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({en_burst_i_34_n_0,en_burst_i_35_n_0,en_burst_i_36_n_0,en_burst_i_37_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_2
       (.CI(en_burst_reg_i_4_n_0),
        .CO({\I_0/en_burst1 ,en_burst_reg_i_2_n_1,en_burst_reg_i_2_n_2,en_burst_reg_i_2_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_burst_i_5_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({en_burst_i_6_n_0,en_burst_i_7_n_0,en_burst_i_8_n_0,en_burst_i_9_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_24
       (.CI(en_burst_reg_i_38_n_0),
        .CO({en_burst_reg_i_24_n_0,en_burst_reg_i_24_n_1,en_burst_reg_i_24_n_2,en_burst_reg_i_24_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_burst_i_39_n_0,en_burst_i_40_n_0,en_burst_i_41_n_0,en_burst_i_42_n_0}),
        .S({en_burst_i_43_n_0,en_burst_i_44_n_0,en_burst_i_45_n_0,en_burst_i_46_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_3
       (.CI(en_burst_reg_i_10_n_0),
        .CO({\I_0/en_burst10_in ,en_burst_reg_i_3_n_1,en_burst_reg_i_3_n_2,en_burst_reg_i_3_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({en_burst_i_11_n_0,en_burst_i_12_n_0,en_burst_i_13_n_0,en_burst_i_14_n_0}),
        .S({en_burst_i_15_n_0,en_burst_i_16_n_0,en_burst_i_17_n_0,en_burst_i_18_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_33
       (.CI(\<const0>__0__0 ),
        .CO({en_burst_reg_i_33_n_0,en_burst_reg_i_33_n_1,en_burst_reg_i_33_n_2,en_burst_reg_i_33_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({en_burst_i_47_n_0,en_burst_i_48_n_0,en_burst_i_49_n_0,en_burst_i_50_n_0}),
        .S({en_burst_i_51_n_0,en_burst_i_52_n_0,en_burst_i_53_n_0,en_burst_i_54_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_38
       (.CI(\<const0>__0__0 ),
        .CO({en_burst_reg_i_38_n_0,en_burst_reg_i_38_n_1,en_burst_reg_i_38_n_2,en_burst_reg_i_38_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({en_burst_i_55_n_0,en_burst_i_56_n_0,en_burst_i_57_n_0,en_burst_i_58_n_0}),
        .S({en_burst_i_59_n_0,en_burst_i_60_n_0,en_burst_i_61_n_0,en_burst_i_62_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 en_burst_reg_i_4
       (.CI(en_burst_reg_i_19_n_0),
        .CO({en_burst_reg_i_4_n_0,en_burst_reg_i_4_n_1,en_burst_reg_i_4_n_2,en_burst_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({en_burst_i_20_n_0,en_burst_i_21_n_0,en_burst_i_22_n_0,en_burst_i_23_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    framereset_i_1
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr0 ),
        .I2(\I_0/i_framereset ),
        .O(framereset_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA954AB54)) 
    g0_b0
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFC666C6660000)) 
    g0_b0__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[3]),
        .I3(in_b[4]),
        .I4(g0_b0_n_0),
        .I5(g0_b0__1_n_0),
        .O(g0_b0__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC66639993999C666)) 
    g0_b0__0__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[3]),
        .I3(in_b[4]),
        .I4(g0_b0__1_n_0),
        .I5(g0_b0_n_0),
        .O(g0_b0__0__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8C6318C6)) 
    g0_b0__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b0__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h64CD9932)) 
    g0_b1
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3C1E1E1E)) 
    g0_b1__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h294A5294)) 
    g0_b1__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h49692DA4)) 
    g0_b2
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA954AB54)) 
    g0_b2__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h318C6318)) 
    g0_b2__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b2__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8E71CE38)) 
    g0_b3
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCE673398)) 
    g0_b3__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h94A5294A)) 
    g0_b3__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b3__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h5AD4A56A)) 
    g0_b4
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0F87C3E0)) 
    g0_b4__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h26C9B26C)) 
    g0_b4__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b4__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6C99364C)) 
    g0_b5
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF007FC00)) 
    g0_b5__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC70E3C70)) 
    g0_b5__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b5__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8F1E3870)) 
    g0_b6
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF80000)) 
    g0_b6__0
       (.I0(in_b[0]),
        .I1(in_b[1]),
        .I2(in_b[2]),
        .I3(in_b[3]),
        .I4(in_b[4]),
        .O(g0_b6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h07F03F80)) 
    g0_b6__1
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b6__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0FE03F80)) 
    g0_b7
       (.I0(in_g[0]),
        .I1(in_g[1]),
        .I2(in_g[2]),
        .I3(in_g[3]),
        .I4(in_g[4]),
        .O(g0_b7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h07FFC000)) 
    g0_b7__0
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3F80)) 
    g0_b8
       (.I0(in_g[1]),
        .I1(in_g[2]),
        .I2(in_g[3]),
        .I3(in_g[4]),
        .O(g0_b8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF8000000)) 
    g0_b8__0
       (.I0(in_r[0]),
        .I1(in_r[1]),
        .I2(in_r[2]),
        .I3(in_r[3]),
        .I4(in_r[4]),
        .O(g0_b8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    g0_b9
       (.I0(in_g[2]),
        .I1(in_g[3]),
        .I2(in_g[4]),
        .O(g0_b9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7F808080)) 
    g0_b9__0
       (.I0(in_g[2]),
        .I1(in_g[3]),
        .I2(in_g[4]),
        .I3(g0_b8__0_n_0),
        .I4(g0_b8_n_0),
        .O(g0_b9__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__0_i_1
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr2_carry__4_n_5 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(hlctr1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__0_i_2
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr2_carry__3_n_4 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(hlctr1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__0_i_3
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr2_carry__3_n_7 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(hlctr1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__0_i_4
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr2_carry__2_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(hlctr1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    hlctr1_carry__1_i_1
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .O(hlctr1_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__1_i_2
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr2_carry__6_n_7 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(hlctr1_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    hlctr1_carry__1_i_3
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr2_carry__5_n_6 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(hlctr1_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    hlctr1_carry_i_1
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr2_carry__1_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(hlctr1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    hlctr1_carry_i_2
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr2_carry__0_n_5 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(hlctr1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    hlctr1_carry_i_3
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(hlctr1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    hlctr1_carry_i_4
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(hlctr1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \hlctr[0]_i_1 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .O(\I_0/hlctr [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[10]_i_1 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[11]_i_1 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[12]_i_1 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[13]_i_1 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[14]_i_1 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[15]_i_1 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[16]_i_1 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[17]_i_1 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[18]_i_1 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[19]_i_1 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[1]_i_1 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[20]_i_1 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[21]_i_1 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[22]_i_1 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[23]_i_1 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[24]_i_1 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[25]_i_1 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[26]_i_1 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[27]_i_1 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[28]_i_1 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[29]_i_1 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[2]_i_1 
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[30]_i_1 
       (.I0(\I_0/hlctr2_carry__6_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55404040)) 
    \hlctr[31]_i_1 
       (.I0(\I_0/i_en_vertbr_last ),
        .I1(\I_0/i_phase4 ),
        .I2(\I_0/i_en_vertbr2 ),
        .I3(\I_0/i_en_vertbr131_in ),
        .I4(\I_0/i_en_vertbr1 ),
        .O(\I_0/hlctr0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[31]_i_2 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[3]_i_1 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[4]_i_1 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[5]_i_1 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[6]_i_1 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[7]_i_1 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[8]_i_1 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \hlctr[9]_i_1 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\I_0/hlctr [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h3A)) 
    i_austastung_i_1
       (.I0(\I_0/i_austastung ),
        .I1(i_austastung_i_3_n_0),
        .I2(\I_0/hlctr0 ),
        .O(i_austastung_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_10
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_austastung_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_11
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_austastung_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_austastung_i_13
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_austastung_i_14
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_austastung_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_15
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_austastung_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_16
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_austastung_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_17
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_austastung_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_19
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_austastung_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    i_austastung_i_2
       (.I0(reset),
        .O(i_austastung_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_20
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_austastung_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_21
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_austastung_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_22
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_austastung_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_24
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_austastung_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_25
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_austastung_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_26
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_austastung_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_27
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_austastung_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_austastung_i_29
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(i_austastung_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000077707770777)) 
    i_austastung_i_3
       (.I0(\I_0/i_sync_c211_in ),
        .I1(\I_0/i_sync_c210_in ),
        .I2(\I_0/i_sync_c2 ),
        .I3(\I_0/i_austastung1 ),
        .I4(\I_0/i_sync_c28_in ),
        .I5(\I_0/i_austastung2 ),
        .O(i_austastung_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_30
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_austastung_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_31
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_austastung_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_32
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_austastung_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_austastung_i_33
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_austastung_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_35
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_austastung_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_36
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_austastung_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_37
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_austastung_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_38
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_austastung_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_austastung_i_39
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_austastung_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_40
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_austastung_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    i_austastung_i_41
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_austastung_i_42
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_5 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_austastung_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_austastung_i_43
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_4 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_austastung_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    i_austastung_i_44
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_austastung_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    i_austastung_i_45
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_austastung_i_46
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_austastung_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    i_austastung_i_47
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_48
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_austastung_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_austastung_i_49
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_austastung_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    i_austastung_i_50
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_austastung_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    i_austastung_i_51
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_austastung_i_7
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_austastung_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_austastung_i_8
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_austastung_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_austastung_i_9
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_austastung_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_12
       (.CI(i_austastung_reg_i_23_n_0),
        .CO({i_austastung_reg_i_12_n_0,i_austastung_reg_i_12_n_1,i_austastung_reg_i_12_n_2,i_austastung_reg_i_12_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_austastung_i_24_n_0,i_austastung_i_25_n_0,i_austastung_i_26_n_0,i_austastung_i_27_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_18
       (.CI(i_austastung_reg_i_28_n_0),
        .CO({i_austastung_reg_i_18_n_0,i_austastung_reg_i_18_n_1,i_austastung_reg_i_18_n_2,i_austastung_reg_i_18_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,i_austastung_i_29_n_0}),
        .S({i_austastung_i_30_n_0,i_austastung_i_31_n_0,i_austastung_i_32_n_0,i_austastung_i_33_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_23
       (.CI(i_austastung_reg_i_34_n_0),
        .CO({i_austastung_reg_i_23_n_0,i_austastung_reg_i_23_n_1,i_austastung_reg_i_23_n_2,i_austastung_reg_i_23_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_austastung_i_35_n_0,i_austastung_i_36_n_0,i_austastung_i_37_n_0,i_austastung_i_38_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_28
       (.CI(\<const0>__0__0 ),
        .CO({i_austastung_reg_i_28_n_0,i_austastung_reg_i_28_n_1,i_austastung_reg_i_28_n_2,i_austastung_reg_i_28_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_austastung_i_39_n_0,i_austastung_i_40_n_0,i_austastung_i_41_n_0,\<const0>__0__0 }),
        .S({i_austastung_i_42_n_0,i_austastung_i_43_n_0,i_austastung_i_44_n_0,i_austastung_i_45_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_34
       (.CI(\<const0>__0__0 ),
        .CO({i_austastung_reg_i_34_n_0,i_austastung_reg_i_34_n_1,i_austastung_reg_i_34_n_2,i_austastung_reg_i_34_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,i_austastung_i_46_n_0,i_austastung_i_47_n_0,\<const0>__0__0 }),
        .S({i_austastung_i_48_n_0,i_austastung_i_49_n_0,i_austastung_i_50_n_0,i_austastung_i_51_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_4
       (.CI(i_austastung_reg_i_6_n_0),
        .CO({\I_0/i_austastung1 ,i_austastung_reg_i_4_n_1,i_austastung_reg_i_4_n_2,i_austastung_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_austastung_i_7_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_austastung_i_8_n_0,i_austastung_i_9_n_0,i_austastung_i_10_n_0,i_austastung_i_11_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_5
       (.CI(i_austastung_reg_i_12_n_0),
        .CO({\I_0/i_austastung2 ,i_austastung_reg_i_5_n_1,i_austastung_reg_i_5_n_2,i_austastung_reg_i_5_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_austastung_i_13_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_austastung_i_14_n_0,i_austastung_i_15_n_0,i_austastung_i_16_n_0,i_austastung_i_17_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_austastung_reg_i_6
       (.CI(i_austastung_reg_i_18_n_0),
        .CO({i_austastung_reg_i_6_n_0,i_austastung_reg_i_6_n_1,i_austastung_reg_i_6_n_2,i_austastung_reg_i_6_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_austastung_i_19_n_0,i_austastung_i_20_n_0,i_austastung_i_21_n_0,i_austastung_i_22_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    i_en_sync_last_i_1
       (.I0(\I_0/i_phase433_in ),
        .I1(\I_0/i_phase4 ),
        .O(\I_0/i_phase3 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_10
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(i_en_sync_last_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_11
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(i_en_sync_last_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_12
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(i_en_sync_last_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_13
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(i_en_sync_last_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_15
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(i_en_sync_last_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_16
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(i_en_sync_last_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_17
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(i_en_sync_last_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_18
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(i_en_sync_last_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_19
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(i_en_sync_last_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_20
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(i_en_sync_last_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_en_sync_last_i_21
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_7 ),
        .O(i_en_sync_last_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    i_en_sync_last_i_22
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(i_en_sync_last_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_23
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(i_en_sync_last_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_sync_last_i_24
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_6 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(i_en_sync_last_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_en_sync_last_i_25
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(i_en_sync_last_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_en_sync_last_i_4
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(i_en_sync_last_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_en_sync_last_i_5
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_en_sync_last_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_6
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(i_en_sync_last_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_7
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(i_en_sync_last_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_sync_last_i_8
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(i_en_sync_last_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_sync_last_reg_i_14
       (.CI(\<const0>__0__0 ),
        .CO({i_en_sync_last_reg_i_14_n_0,i_en_sync_last_reg_i_14_n_1,i_en_sync_last_reg_i_14_n_2,i_en_sync_last_reg_i_14_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_en_sync_last_i_19_n_0,\<const0>__0__0 ,i_en_sync_last_i_20_n_0,i_en_sync_last_i_21_n_0}),
        .S({i_en_sync_last_i_22_n_0,i_en_sync_last_i_23_n_0,i_en_sync_last_i_24_n_0,i_en_sync_last_i_25_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_sync_last_reg_i_2
       (.CI(i_en_sync_last_reg_i_3_n_0),
        .CO({\I_0/i_phase433_in ,i_en_sync_last_reg_i_2_n_1,i_en_sync_last_reg_i_2_n_2,i_en_sync_last_reg_i_2_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_sync_last_i_4_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_sync_last_i_5_n_0,i_en_sync_last_i_6_n_0,i_en_sync_last_i_7_n_0,i_en_sync_last_i_8_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_sync_last_reg_i_3
       (.CI(i_en_sync_last_reg_i_9_n_0),
        .CO({i_en_sync_last_reg_i_3_n_0,i_en_sync_last_reg_i_3_n_1,i_en_sync_last_reg_i_3_n_2,i_en_sync_last_reg_i_3_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_sync_last_i_10_n_0,i_en_sync_last_i_11_n_0,i_en_sync_last_i_12_n_0,i_en_sync_last_i_13_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_sync_last_reg_i_9
       (.CI(i_en_sync_last_reg_i_14_n_0),
        .CO({i_en_sync_last_reg_i_9_n_0,i_en_sync_last_reg_i_9_n_1,i_en_sync_last_reg_i_9_n_2,i_en_sync_last_reg_i_9_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_sync_last_i_15_n_0,i_en_sync_last_i_16_n_0,i_en_sync_last_i_17_n_0,i_en_sync_last_i_18_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    i_en_vertbr_last_i_1
       (.I0(\I_0/i_phase4 ),
        .I1(\I_0/i_en_vertbr2 ),
        .I2(\I_0/i_en_vertbr131_in ),
        .I3(\I_0/i_en_vertbr1 ),
        .O(\I_0/i_en_vertbr ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_10
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(i_en_vertbr_last_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_en_vertbr_last_i_12
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(i_en_vertbr_last_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_en_vertbr_last_i_13
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_en_vertbr_last_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_14
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(i_en_vertbr_last_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_15
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(i_en_vertbr_last_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_16
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(i_en_vertbr_last_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_18
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_en_vertbr_last_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_19
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__6_n_7 ),
        .O(i_en_vertbr_last_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_20
       (.I0(\I_0/pixctr2_carry__5_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_5 ),
        .O(i_en_vertbr_last_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_21
       (.I0(\I_0/pixctr2_carry__4_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_7 ),
        .O(i_en_vertbr_last_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_en_vertbr_last_i_22
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_en_vertbr_last_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_23
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(i_en_vertbr_last_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_24
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(i_en_vertbr_last_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_25
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(i_en_vertbr_last_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_27
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(i_en_vertbr_last_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_28
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(i_en_vertbr_last_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_29
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(i_en_vertbr_last_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_30
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(i_en_vertbr_last_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_32
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(i_en_vertbr_last_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_33
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(i_en_vertbr_last_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_34
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(i_en_vertbr_last_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_35
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(i_en_vertbr_last_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_37
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_5 ),
        .O(i_en_vertbr_last_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_38
       (.I0(\I_0/pixctr2_carry__3_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_7 ),
        .O(i_en_vertbr_last_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_39
       (.I0(\I_0/pixctr2_carry__3_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_5 ),
        .O(i_en_vertbr_last_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_40
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_7 ),
        .O(i_en_vertbr_last_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_41
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(i_en_vertbr_last_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_42
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(i_en_vertbr_last_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_43
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(i_en_vertbr_last_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_44
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(i_en_vertbr_last_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_46
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(i_en_vertbr_last_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_47
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(i_en_vertbr_last_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_48
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(i_en_vertbr_last_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_49
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(i_en_vertbr_last_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_50
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(i_en_vertbr_last_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    i_en_vertbr_last_i_52
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr1_carry__1_n_1 ),
        .O(i_en_vertbr_last_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_53
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(i_en_vertbr_last_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_54
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(i_en_vertbr_last_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_55
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(i_en_vertbr_last_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    i_en_vertbr_last_i_56
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(i_en_vertbr_last_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_58
       (.I0(\I_0/pixctr2_carry__2_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_5 ),
        .O(i_en_vertbr_last_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_59
       (.I0(\I_0/pixctr2_carry__1_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_7 ),
        .O(i_en_vertbr_last_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_en_vertbr_last_i_6
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(i_en_vertbr_last_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_60
       (.I0(\I_0/pixctr2_carry__1_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_5 ),
        .O(i_en_vertbr_last_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_en_vertbr_last_i_61
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(i_en_vertbr_last_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_62
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(i_en_vertbr_last_i_62_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_63
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(i_en_vertbr_last_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_64
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(i_en_vertbr_last_i_64_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_65
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_4 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(i_en_vertbr_last_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_en_vertbr_last_i_66
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .O(i_en_vertbr_last_i_66_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_67
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(i_en_vertbr_last_i_67_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_en_vertbr_last_i_68
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .O(i_en_vertbr_last_i_68_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_69
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(i_en_vertbr_last_i_69_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_en_vertbr_last_i_7
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_en_vertbr_last_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    i_en_vertbr_last_i_70
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(i_en_vertbr_last_i_70_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_71
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(i_en_vertbr_last_i_71_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCE)) 
    i_en_vertbr_last_i_72
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(i_en_vertbr_last_i_72_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_73
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(i_en_vertbr_last_i_73_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    i_en_vertbr_last_i_74
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(i_en_vertbr_last_i_74_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_en_vertbr_last_i_75
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .O(i_en_vertbr_last_i_75_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    i_en_vertbr_last_i_76
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(i_en_vertbr_last_i_76_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_en_vertbr_last_i_77
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(i_en_vertbr_last_i_77_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_78
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_5 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(i_en_vertbr_last_i_78_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCE)) 
    i_en_vertbr_last_i_79
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(i_en_vertbr_last_i_79_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_8
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(i_en_vertbr_last_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_en_vertbr_last_i_80
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(i_en_vertbr_last_i_80_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_en_vertbr_last_i_81
       (.I0(\I_0/pixctr2_carry_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(i_en_vertbr_last_i_81_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h23)) 
    i_en_vertbr_last_i_82
       (.I0(\I_0/pixctr2_carry_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr_reg_n_0_ ),
        .O(i_en_vertbr_last_i_82_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_en_vertbr_last_i_83
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(i_en_vertbr_last_i_83_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_en_vertbr_last_i_84
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(i_en_vertbr_last_i_84_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_85
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(i_en_vertbr_last_i_85_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCE)) 
    i_en_vertbr_last_i_86
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(i_en_vertbr_last_i_86_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_en_vertbr_last_i_9
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(i_en_vertbr_last_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_11
       (.CI(i_en_vertbr_last_reg_i_31_n_0),
        .CO({i_en_vertbr_last_reg_i_11_n_0,i_en_vertbr_last_reg_i_11_n_1,i_en_vertbr_last_reg_i_11_n_2,i_en_vertbr_last_reg_i_11_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_32_n_0,i_en_vertbr_last_i_33_n_0,i_en_vertbr_last_i_34_n_0,i_en_vertbr_last_i_35_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_17
       (.CI(i_en_vertbr_last_reg_i_36_n_0),
        .CO({i_en_vertbr_last_reg_i_17_n_0,i_en_vertbr_last_reg_i_17_n_1,i_en_vertbr_last_reg_i_17_n_2,i_en_vertbr_last_reg_i_17_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_vertbr_last_i_37_n_0,i_en_vertbr_last_i_38_n_0,i_en_vertbr_last_i_39_n_0,i_en_vertbr_last_i_40_n_0}),
        .S({i_en_vertbr_last_i_41_n_0,i_en_vertbr_last_i_42_n_0,i_en_vertbr_last_i_43_n_0,i_en_vertbr_last_i_44_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_2
       (.CI(i_en_vertbr_last_reg_i_5_n_0),
        .CO({\I_0/i_en_vertbr2 ,i_en_vertbr_last_reg_i_2_n_1,i_en_vertbr_last_reg_i_2_n_2,i_en_vertbr_last_reg_i_2_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_vertbr_last_i_6_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_7_n_0,i_en_vertbr_last_i_8_n_0,i_en_vertbr_last_i_9_n_0,i_en_vertbr_last_i_10_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_26
       (.CI(i_en_vertbr_last_reg_i_45_n_0),
        .CO({i_en_vertbr_last_reg_i_26_n_0,i_en_vertbr_last_reg_i_26_n_1,i_en_vertbr_last_reg_i_26_n_2,i_en_vertbr_last_reg_i_26_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,i_en_vertbr_last_i_46_n_0}),
        .S({i_en_vertbr_last_i_47_n_0,i_en_vertbr_last_i_48_n_0,i_en_vertbr_last_i_49_n_0,i_en_vertbr_last_i_50_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_3
       (.CI(i_en_vertbr_last_reg_i_11_n_0),
        .CO({\I_0/i_en_vertbr131_in ,i_en_vertbr_last_reg_i_3_n_1,i_en_vertbr_last_reg_i_3_n_2,i_en_vertbr_last_reg_i_3_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_vertbr_last_i_12_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_13_n_0,i_en_vertbr_last_i_14_n_0,i_en_vertbr_last_i_15_n_0,i_en_vertbr_last_i_16_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_31
       (.CI(i_en_vertbr_last_reg_i_51_n_0),
        .CO({i_en_vertbr_last_reg_i_31_n_0,i_en_vertbr_last_reg_i_31_n_1,i_en_vertbr_last_reg_i_31_n_2,i_en_vertbr_last_reg_i_31_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,i_en_vertbr_last_i_52_n_0}),
        .S({i_en_vertbr_last_i_53_n_0,i_en_vertbr_last_i_54_n_0,i_en_vertbr_last_i_55_n_0,i_en_vertbr_last_i_56_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_36
       (.CI(i_en_vertbr_last_reg_i_57_n_0),
        .CO({i_en_vertbr_last_reg_i_36_n_0,i_en_vertbr_last_reg_i_36_n_1,i_en_vertbr_last_reg_i_36_n_2,i_en_vertbr_last_reg_i_36_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_vertbr_last_i_58_n_0,i_en_vertbr_last_i_59_n_0,i_en_vertbr_last_i_60_n_0,i_en_vertbr_last_i_61_n_0}),
        .S({i_en_vertbr_last_i_62_n_0,i_en_vertbr_last_i_63_n_0,i_en_vertbr_last_i_64_n_0,i_en_vertbr_last_i_65_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_4
       (.CI(i_en_vertbr_last_reg_i_17_n_0),
        .CO({\I_0/i_en_vertbr1 ,i_en_vertbr_last_reg_i_4_n_1,i_en_vertbr_last_reg_i_4_n_2,i_en_vertbr_last_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_en_vertbr_last_i_18_n_0,i_en_vertbr_last_i_19_n_0,i_en_vertbr_last_i_20_n_0,i_en_vertbr_last_i_21_n_0}),
        .S({i_en_vertbr_last_i_22_n_0,i_en_vertbr_last_i_23_n_0,i_en_vertbr_last_i_24_n_0,i_en_vertbr_last_i_25_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_45
       (.CI(\<const0>__0__0 ),
        .CO({i_en_vertbr_last_reg_i_45_n_0,i_en_vertbr_last_reg_i_45_n_1,i_en_vertbr_last_reg_i_45_n_2,i_en_vertbr_last_reg_i_45_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_en_vertbr_last_i_66_n_0,i_en_vertbr_last_i_67_n_0,i_en_vertbr_last_i_68_n_0,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_69_n_0,i_en_vertbr_last_i_70_n_0,i_en_vertbr_last_i_71_n_0,i_en_vertbr_last_i_72_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_5
       (.CI(i_en_vertbr_last_reg_i_26_n_0),
        .CO({i_en_vertbr_last_reg_i_5_n_0,i_en_vertbr_last_reg_i_5_n_1,i_en_vertbr_last_reg_i_5_n_2,i_en_vertbr_last_reg_i_5_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_27_n_0,i_en_vertbr_last_i_28_n_0,i_en_vertbr_last_i_29_n_0,i_en_vertbr_last_i_30_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_51
       (.CI(\<const0>__0__0 ),
        .CO({i_en_vertbr_last_reg_i_51_n_0,i_en_vertbr_last_reg_i_51_n_1,i_en_vertbr_last_reg_i_51_n_2,i_en_vertbr_last_reg_i_51_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_en_vertbr_last_i_73_n_0,i_en_vertbr_last_i_74_n_0,i_en_vertbr_last_i_75_n_0,\<const0>__0__0 }),
        .S({i_en_vertbr_last_i_76_n_0,i_en_vertbr_last_i_77_n_0,i_en_vertbr_last_i_78_n_0,i_en_vertbr_last_i_79_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_en_vertbr_last_reg_i_57
       (.CI(\<const0>__0__0 ),
        .CO({i_en_vertbr_last_reg_i_57_n_0,i_en_vertbr_last_reg_i_57_n_1,i_en_vertbr_last_reg_i_57_n_2,i_en_vertbr_last_reg_i_57_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,i_en_vertbr_last_i_80_n_0,i_en_vertbr_last_i_81_n_0,i_en_vertbr_last_i_82_n_0}),
        .S({i_en_vertbr_last_i_83_n_0,i_en_vertbr_last_i_84_n_0,i_en_vertbr_last_i_85_n_0,i_en_vertbr_last_i_86_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__0_i_1
       (.I0(\I_0/pixctr2_carry__2_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_5 ),
        .O(i_phase4_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__0_i_2
       (.I0(\I_0/pixctr2_carry__1_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_7 ),
        .O(i_phase4_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__0_i_3
       (.I0(\I_0/pixctr2_carry__1_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_5 ),
        .O(i_phase4_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__0_i_4
       (.I0(\I_0/pixctr2_carry__0_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_7 ),
        .O(i_phase4_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__0_i_5
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(i_phase4_inferred__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__0_i_6
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(i_phase4_inferred__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__0_i_7
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(i_phase4_inferred__0_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__0_i_8
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(i_phase4_inferred__0_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__1_i_1
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_5 ),
        .O(i_phase4_inferred__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__1_i_2
       (.I0(\I_0/pixctr2_carry__3_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_7 ),
        .O(i_phase4_inferred__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__1_i_3
       (.I0(\I_0/pixctr2_carry__3_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_5 ),
        .O(i_phase4_inferred__0_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__1_i_4
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_7 ),
        .O(i_phase4_inferred__0_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__1_i_5
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(i_phase4_inferred__0_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__1_i_6
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(i_phase4_inferred__0_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__1_i_7
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(i_phase4_inferred__0_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__1_i_8
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(i_phase4_inferred__0_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_phase4_inferred__0_carry__2_i_1
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_phase4_inferred__0_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__2_i_2
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__6_n_7 ),
        .O(i_phase4_inferred__0_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__2_i_3
       (.I0(\I_0/pixctr2_carry__5_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_5 ),
        .O(i_phase4_inferred__0_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry__2_i_4
       (.I0(\I_0/pixctr2_carry__4_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_7 ),
        .O(i_phase4_inferred__0_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_phase4_inferred__0_carry__2_i_5
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(i_phase4_inferred__0_carry__2_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__2_i_6
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(i_phase4_inferred__0_carry__2_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__2_i_7
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(i_phase4_inferred__0_carry__2_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry__2_i_8
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(i_phase4_inferred__0_carry__2_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry_i_1
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_5 ),
        .O(i_phase4_inferred__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry_i_2
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_7 ),
        .O(i_phase4_inferred__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_phase4_inferred__0_carry_i_3
       (.I0(\I_0/pixctr2_carry_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(i_phase4_inferred__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h23)) 
    i_phase4_inferred__0_carry_i_4
       (.I0(\I_0/pixctr2_carry_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr_reg_n_0_ ),
        .O(i_phase4_inferred__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry_i_5
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(i_phase4_inferred__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry_i_6
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(i_phase4_inferred__0_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_phase4_inferred__0_carry_i_7
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(i_phase4_inferred__0_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCE)) 
    i_phase4_inferred__0_carry_i_8
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(i_phase4_inferred__0_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h95AA)) 
    i_phase_i_1
       (.I0(phase),
        .I1(\I_0/i_phase433_in ),
        .I2(\I_0/i_phase4 ),
        .I3(\I_0/i_en_sync_last ),
        .O(i_phase_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    i_phase_i_2
       (.I0(reset),
        .O(i_phase_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF888FFFFF8880000)) 
    i_readmem_i_1
       (.I0(\I_0/i_readmem15_in ),
        .I1(\I_0/i_readmem1 ),
        .I2(\I_0/i_readmem26_in ),
        .I3(\I_0/i_readmem2 ),
        .I4(\I_0/hlctr0 ),
        .I5(readmem),
        .O(i_readmem_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_10
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(i_readmem_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    i_readmem_i_100
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_100_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    i_readmem_i_101
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_readmem_i_101_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_102
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_readmem_i_102_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_readmem_i_103
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .O(i_readmem_i_103_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    i_readmem_i_104
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_104_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_readmem_i_105
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_readmem_i_105_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_106
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_4 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_readmem_i_106_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_107
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_readmem_i_107_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    i_readmem_i_108
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(i_readmem_i_108_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_109
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_readmem_i_109_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_readmem_i_11
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_readmem_i_110
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_readmem_i_110_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    i_readmem_i_111
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_readmem_i_111_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_112
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(i_readmem_i_112_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_113
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_readmem_i_113_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_114
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_readmem_i_114_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_115
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_readmem_i_115_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    i_readmem_i_116
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_116_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_117
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_readmem_i_117_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_readmem_i_118
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_readmem_i_118_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_readmem_i_119
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .O(i_readmem_i_119_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_12
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_readmem_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    i_readmem_i_120
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_120_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_121
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_readmem_i_121_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_122
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_readmem_i_122_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_123
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_readmem_i_123_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    i_readmem_i_124
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(i_readmem_i_124_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_13
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_readmem_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_14
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_readmem_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_readmem_i_16
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_readmem_i_17
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_18
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_readmem_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_19
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_readmem_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_20
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_readmem_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_22
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_23
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(i_readmem_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_24
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(i_readmem_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_25
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(i_readmem_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_readmem_i_26
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_27
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_readmem_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_28
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_readmem_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_29
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_readmem_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_readmem_i_31
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_readmem_i_32
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_33
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_readmem_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_34
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_readmem_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_35
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_readmem_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_37
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(i_readmem_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_38
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(i_readmem_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_39
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(i_readmem_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_40
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(i_readmem_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_41
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_readmem_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_42
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_readmem_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_43
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_readmem_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_44
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_readmem_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_46
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_readmem_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_47
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_readmem_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_48
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_readmem_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_49
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_readmem_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_51
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(i_readmem_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_52
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(i_readmem_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_53
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(i_readmem_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_54
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(i_readmem_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_55
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_readmem_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_56
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_readmem_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_57
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_readmem_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_58
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_readmem_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_60
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_readmem_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_61
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_readmem_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_62
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_readmem_i_62_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_63
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_readmem_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_65
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(i_readmem_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_66
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(i_readmem_i_66_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_67
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(i_readmem_i_67_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_readmem_i_68
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(i_readmem_i_68_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_69
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_readmem_i_69_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_7
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_readmem_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_70
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_readmem_i_70_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_71
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_readmem_i_71_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_72
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_readmem_i_72_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_74
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_readmem_i_74_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_75
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_readmem_i_75_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_76
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_readmem_i_76_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_77
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(i_readmem_i_77_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_78
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_readmem_i_78_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_8
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(i_readmem_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_80
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(i_readmem_i_80_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_81
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(i_readmem_i_81_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_82
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(i_readmem_i_82_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_83
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(i_readmem_i_83_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_84
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_readmem_i_84_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_85
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_readmem_i_85_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_86
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_readmem_i_86_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_87
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_readmem_i_87_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_readmem_i_89
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(i_readmem_i_89_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    i_readmem_i_9
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(i_readmem_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_90
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_readmem_i_90_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_91
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_readmem_i_91_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_readmem_i_92
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_readmem_i_92_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_93
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_readmem_i_93_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    i_readmem_i_94
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_readmem_i_94_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_readmem_i_95
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_readmem_i_95_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h51)) 
    i_readmem_i_96
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(i_readmem_i_96_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_97
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_5 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_readmem_i_97_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_readmem_i_98
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_4 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_readmem_i_98_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    i_readmem_i_99
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_readmem_i_99_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_15
       (.CI(i_readmem_reg_i_45_n_0),
        .CO({i_readmem_reg_i_15_n_0,i_readmem_reg_i_15_n_1,i_readmem_reg_i_15_n_2,i_readmem_reg_i_15_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_readmem_i_46_n_0,i_readmem_i_47_n_0,i_readmem_i_48_n_0,i_readmem_i_49_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_2
       (.CI(i_readmem_reg_i_6_n_0),
        .CO({\I_0/i_readmem15_in ,i_readmem_reg_i_2_n_1,i_readmem_reg_i_2_n_2,i_readmem_reg_i_2_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_7_n_0,i_readmem_i_8_n_0,i_readmem_i_9_n_0,i_readmem_i_10_n_0}),
        .S({i_readmem_i_11_n_0,i_readmem_i_12_n_0,i_readmem_i_13_n_0,i_readmem_i_14_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_21
       (.CI(i_readmem_reg_i_50_n_0),
        .CO({i_readmem_reg_i_21_n_0,i_readmem_reg_i_21_n_1,i_readmem_reg_i_21_n_2,i_readmem_reg_i_21_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_51_n_0,i_readmem_i_52_n_0,i_readmem_i_53_n_0,i_readmem_i_54_n_0}),
        .S({i_readmem_i_55_n_0,i_readmem_i_56_n_0,i_readmem_i_57_n_0,i_readmem_i_58_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_3
       (.CI(i_readmem_reg_i_15_n_0),
        .CO({\I_0/i_readmem1 ,i_readmem_reg_i_3_n_1,i_readmem_reg_i_3_n_2,i_readmem_reg_i_3_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_16_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_readmem_i_17_n_0,i_readmem_i_18_n_0,i_readmem_i_19_n_0,i_readmem_i_20_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_30
       (.CI(i_readmem_reg_i_59_n_0),
        .CO({i_readmem_reg_i_30_n_0,i_readmem_reg_i_30_n_1,i_readmem_reg_i_30_n_2,i_readmem_reg_i_30_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_readmem_i_60_n_0,i_readmem_i_61_n_0,i_readmem_i_62_n_0,i_readmem_i_63_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_36
       (.CI(i_readmem_reg_i_64_n_0),
        .CO({i_readmem_reg_i_36_n_0,i_readmem_reg_i_36_n_1,i_readmem_reg_i_36_n_2,i_readmem_reg_i_36_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_65_n_0,i_readmem_i_66_n_0,i_readmem_i_67_n_0,i_readmem_i_68_n_0}),
        .S({i_readmem_i_69_n_0,i_readmem_i_70_n_0,i_readmem_i_71_n_0,i_readmem_i_72_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_4
       (.CI(i_readmem_reg_i_21_n_0),
        .CO({\I_0/i_readmem26_in ,i_readmem_reg_i_4_n_1,i_readmem_reg_i_4_n_2,i_readmem_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_22_n_0,i_readmem_i_23_n_0,i_readmem_i_24_n_0,i_readmem_i_25_n_0}),
        .S({i_readmem_i_26_n_0,i_readmem_i_27_n_0,i_readmem_i_28_n_0,i_readmem_i_29_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_45
       (.CI(i_readmem_reg_i_73_n_0),
        .CO({i_readmem_reg_i_45_n_0,i_readmem_reg_i_45_n_1,i_readmem_reg_i_45_n_2,i_readmem_reg_i_45_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,i_readmem_i_74_n_0,\<const0>__0__0 }),
        .S({i_readmem_i_75_n_0,i_readmem_i_76_n_0,i_readmem_i_77_n_0,i_readmem_i_78_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_5
       (.CI(i_readmem_reg_i_30_n_0),
        .CO({\I_0/i_readmem2 ,i_readmem_reg_i_5_n_1,i_readmem_reg_i_5_n_2,i_readmem_reg_i_5_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_31_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({i_readmem_i_32_n_0,i_readmem_i_33_n_0,i_readmem_i_34_n_0,i_readmem_i_35_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_50
       (.CI(i_readmem_reg_i_79_n_0),
        .CO({i_readmem_reg_i_50_n_0,i_readmem_reg_i_50_n_1,i_readmem_reg_i_50_n_2,i_readmem_reg_i_50_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_80_n_0,i_readmem_i_81_n_0,i_readmem_i_82_n_0,i_readmem_i_83_n_0}),
        .S({i_readmem_i_84_n_0,i_readmem_i_85_n_0,i_readmem_i_86_n_0,i_readmem_i_87_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_59
       (.CI(i_readmem_reg_i_88_n_0),
        .CO({i_readmem_reg_i_59_n_0,i_readmem_reg_i_59_n_1,i_readmem_reg_i_59_n_2,i_readmem_reg_i_59_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,i_readmem_i_89_n_0}),
        .S({i_readmem_i_90_n_0,i_readmem_i_91_n_0,i_readmem_i_92_n_0,i_readmem_i_93_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_6
       (.CI(i_readmem_reg_i_36_n_0),
        .CO({i_readmem_reg_i_6_n_0,i_readmem_reg_i_6_n_1,i_readmem_reg_i_6_n_2,i_readmem_reg_i_6_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({i_readmem_i_37_n_0,i_readmem_i_38_n_0,i_readmem_i_39_n_0,i_readmem_i_40_n_0}),
        .S({i_readmem_i_41_n_0,i_readmem_i_42_n_0,i_readmem_i_43_n_0,i_readmem_i_44_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_64
       (.CI(\<const0>__0__0 ),
        .CO({i_readmem_reg_i_64_n_0,i_readmem_reg_i_64_n_1,i_readmem_reg_i_64_n_2,i_readmem_reg_i_64_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_readmem_i_94_n_0,i_readmem_i_95_n_0,\<const0>__0__0 ,i_readmem_i_96_n_0}),
        .S({i_readmem_i_97_n_0,i_readmem_i_98_n_0,i_readmem_i_99_n_0,i_readmem_i_100_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_73
       (.CI(\<const0>__0__0 ),
        .CO({i_readmem_reg_i_73_n_0,i_readmem_reg_i_73_n_1,i_readmem_reg_i_73_n_2,i_readmem_reg_i_73_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_readmem_i_101_n_0,i_readmem_i_102_n_0,i_readmem_i_103_n_0,i_readmem_i_104_n_0}),
        .S({i_readmem_i_105_n_0,i_readmem_i_106_n_0,i_readmem_i_107_n_0,i_readmem_i_108_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_79
       (.CI(\<const0>__0__0 ),
        .CO({i_readmem_reg_i_79_n_0,i_readmem_reg_i_79_n_1,i_readmem_reg_i_79_n_2,i_readmem_reg_i_79_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_readmem_i_109_n_0,i_readmem_i_110_n_0,i_readmem_i_111_n_0,i_readmem_i_112_n_0}),
        .S({i_readmem_i_113_n_0,i_readmem_i_114_n_0,i_readmem_i_115_n_0,i_readmem_i_116_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 i_readmem_reg_i_88
       (.CI(\<const0>__0__0 ),
        .CO({i_readmem_reg_i_88_n_0,i_readmem_reg_i_88_n_1,i_readmem_reg_i_88_n_2,i_readmem_reg_i_88_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({i_readmem_i_117_n_0,i_readmem_i_118_n_0,i_readmem_i_119_n_0,i_readmem_i_120_n_0}),
        .S({i_readmem_i_121_n_0,i_readmem_i_122_n_0,i_readmem_i_123_n_0,i_readmem_i_124_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_sync_c2_inferred__9_carry__0_i_1
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(i_sync_c2_inferred__9_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__0_i_2
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(i_sync_c2_inferred__9_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__0_i_3
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(i_sync_c2_inferred__9_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__0_i_4
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(i_sync_c2_inferred__9_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_sync_c2_inferred__9_carry__0_i_5
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(i_sync_c2_inferred__9_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__1_i_1
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(i_sync_c2_inferred__9_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__1_i_2
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(i_sync_c2_inferred__9_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__1_i_3
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(i_sync_c2_inferred__9_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__1_i_4
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(i_sync_c2_inferred__9_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    i_sync_c2_inferred__9_carry__2_i_1
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_sync_c2_inferred__9_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    i_sync_c2_inferred__9_carry__2_i_2
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(i_sync_c2_inferred__9_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__2_i_3
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(i_sync_c2_inferred__9_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__2_i_4
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(i_sync_c2_inferred__9_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry__2_i_5
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(i_sync_c2_inferred__9_carry__2_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    i_sync_c2_inferred__9_carry_i_1
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(i_sync_c2_inferred__9_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_sync_c2_inferred__9_carry_i_2
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .O(i_sync_c2_inferred__9_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    i_sync_c2_inferred__9_carry_i_3
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .O(i_sync_c2_inferred__9_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    i_sync_c2_inferred__9_carry_i_4
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(i_sync_c2_inferred__9_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_sync_c2_inferred__9_carry_i_5
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(i_sync_c2_inferred__9_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_sync_c2_inferred__9_carry_i_6
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(i_sync_c2_inferred__9_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_sync_c2_inferred__9_carry_i_7
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(i_sync_c2_inferred__9_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    i_sync_c2_inferred__9_carry_i_8
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(i_sync_c2_inferred__9_carry_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8FFF8F00)) 
    \i_sync_c[0]_i_1 
       (.I0(\i_sync_c[0]_i_2_n_0 ),
        .I1(\i_sync_c[0]_i_3_n_0 ),
        .I2(\i_sync_c[0]_i_4_n_0 ),
        .I3(\I_0/hlctr0 ),
        .I4(\I_0/i_sync_c [0]),
        .O(i_sync_c));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF088808880888)) 
    \i_sync_c[0]_i_2 
       (.I0(\I_0/i_sync_c212_in ),
        .I1(\I_0/i_sync_c213_in ),
        .I2(\I_0/i_sync_c215_in ),
        .I3(\I_0/i_sync_c216_in ),
        .I4(\I_0/i_sync_c219_in ),
        .I5(\I_0/i_sync_c218_in ),
        .O(\i_sync_c[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0777)) 
    \i_sync_c[0]_i_3 
       (.I0(\I_0/i_sync_c2 ),
        .I1(\I_0/i_sync_c221_in ),
        .I2(\I_0/i_sync_c227_in ),
        .I3(\I_0/i_sync_c226_in ),
        .O(\i_sync_c[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000F777F777F777)) 
    \i_sync_c[0]_i_4 
       (.I0(\I_0/i_sync_c223_in ),
        .I1(\I_0/i_sync_c224_in ),
        .I2(\I_0/i_sync_c226_in ),
        .I3(\I_0/i_sync_c227_in ),
        .I4(\I_0/i_sync_c28_in ),
        .I5(\I_0/i_sync_c229_in ),
        .O(\i_sync_c[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00750075FFFF0000)) 
    \i_sync_c[1]_i_1 
       (.I0(\i_sync_c[1]_i_2_n_0 ),
        .I1(\i_sync_c[1]_i_3_n_0 ),
        .I2(\i_sync_c[1]_i_4_n_0 ),
        .I3(\i_sync_c[1]_i_5_n_0 ),
        .I4(\I_0/i_sync_c [1]),
        .I5(\I_0/hlctr0 ),
        .O(\i_sync_c[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_100 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_101 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_102 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_103 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_104 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_106 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_107 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_108 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_109 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_110 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_112 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_113 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_114 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_115 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_116 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_117 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_118 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_119 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_119_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_121 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_121_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_122 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_122_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_123 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_123_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_124 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_124_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_125 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_125_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_127 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_127_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_128 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_128_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_129 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_129_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_130 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_130_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_131 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_131_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_132 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_132_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_133 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_133_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_134 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_134_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_136 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_136_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_137 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_137_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_138 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_138_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_139 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_139_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_141 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_142 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_143 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_144 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_145 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_145_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_146 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_146_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_147 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_147_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_148 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_148_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_150 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_150_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_151 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_151_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_152 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_152_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_153 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_153_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_155 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_155_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_156 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_156_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_157 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_157_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_158 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_158_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_159 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_159_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_160 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_160_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_161 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_161_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_162 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_162_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_164 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_164_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_165 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_165_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_166 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_166_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_167 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_167_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_168 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_168_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_169 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_169_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_170 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_170_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_171 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_171_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_173 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_173_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_174 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_174_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_175 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_175_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_176 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_176_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_177 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_177_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_178 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_178_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_179 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_179_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_180 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_180_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_182 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_182_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_183 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_183_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_184 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_184_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_185 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_185_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_187 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_187_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_188 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_188_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_189 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_189_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_190 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_190_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_192 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_192_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_193 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_193_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_194 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_194_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_195 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_195_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_196 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_196_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_197 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_197_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_198 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_198_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_199 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_199_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000077707770777)) 
    \i_sync_c[1]_i_2 
       (.I0(\I_0/i_sync_c226_in ),
        .I1(\I_0/i_sync_c227_in ),
        .I2(\I_0/i_sync_c221_in ),
        .I3(\I_0/i_sync_c2 ),
        .I4(\I_0/i_sync_c224_in ),
        .I5(\I_0/i_sync_c223_in ),
        .O(\i_sync_c[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_201 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_201_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_202 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_202_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_203 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_203_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_204 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_204_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_206 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_206_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_207 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_207_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_208 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_208_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_209 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_209_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_210 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_210_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_211 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_211_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_212 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_212_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_213 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_213_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_215 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_215_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_216 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_216_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_217 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_217_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_218 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_218_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_22 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_220 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_220_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_221 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_221_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_222 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_222_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_223 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_223_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_224 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_224_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_225 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_225_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_226 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_226_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_227 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_227_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_229 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_229_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_23 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_230 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_230_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_231 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_231_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_232 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_232_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_234 
       (.I0(\I_0/hlctr2_carry__4_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_5 ),
        .O(\i_sync_c[1]_i_234_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_235 
       (.I0(\I_0/hlctr2_carry__3_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_7 ),
        .O(\i_sync_c[1]_i_235_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_236 
       (.I0(\I_0/hlctr2_carry__3_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_5 ),
        .O(\i_sync_c[1]_i_236_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_237 
       (.I0(\I_0/hlctr2_carry__2_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_7 ),
        .O(\i_sync_c[1]_i_237_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_238 
       (.I0(\I_0/hlctr2_carry__4_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_6 ),
        .O(\i_sync_c[1]_i_238_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_239 
       (.I0(\I_0/hlctr2_carry__4_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_4 ),
        .O(\i_sync_c[1]_i_239_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_24 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_240 
       (.I0(\I_0/hlctr2_carry__3_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__3_n_6 ),
        .O(\i_sync_c[1]_i_240_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_241 
       (.I0(\I_0/hlctr2_carry__3_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_4 ),
        .O(\i_sync_c[1]_i_241_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_243 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_243_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_244 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_244_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_245 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_245_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_246 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_246_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_248 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_248_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_249 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_249_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_25 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_250 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_250_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_251 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_251_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_252 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_252_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_253 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_253_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_254 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_254_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_255 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_255_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_257 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_257_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_258 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_258_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_259 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_259_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_26 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_260 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_260_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_261 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_261_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_263 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_263_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_264 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_264_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_265 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_265_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_266 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_266_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_267 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_267_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_268 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_268_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_269 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_269_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_270 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_270_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_272 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_272_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_273 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_273_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_274 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_274_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_275 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_275_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_276 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_276_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_277 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_277_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_278 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_278_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_279 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_279_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_28 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_281 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_281_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_282 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_282_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_283 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_283_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_284 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_284_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_285 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_285_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_286 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_286_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_287 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_287_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_288 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_288_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_29 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_290 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_290_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_291 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_291_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_292 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_292_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_293 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_293_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_294 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_294_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_296 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_296_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_297 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_297_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_298 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_298_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_299 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_299_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000077707770777)) 
    \i_sync_c[1]_i_3 
       (.I0(\I_0/i_sync_c213_in ),
        .I1(\I_0/i_sync_c212_in ),
        .I2(\I_0/i_sync_c210_in ),
        .I3(\I_0/i_sync_c211_in ),
        .I4(\I_0/i_sync_c215_in ),
        .I5(\I_0/i_sync_c216_in ),
        .O(\i_sync_c[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_30 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_300 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_300_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_302 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_302_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_303 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_303_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_304 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_304_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_305 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_305_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_306 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_306_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_307 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_307_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_308 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_6 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_308_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_309 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_309_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_31 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_311 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_311_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_312 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_312_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_313 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_313_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_314 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_314_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_315 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_315_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_317 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_317_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_318 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_318_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_319 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_319_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_32 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_320 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_320_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_321 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_321_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_322 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_322_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_323 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_323_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_324 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_324_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_326 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_326_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_327 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_327_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_328 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_328_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_329 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_329_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_33 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_330 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_330_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_332 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_332_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_333 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_333_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_334 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_334_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_335 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_335_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_336 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_336_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_337 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_337_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_338 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_338_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_339 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__1_n_7 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_339_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_34 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_341 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_341_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_342 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_342_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_343 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_343_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_344 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_344_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_346 
       (.I0(\I_0/hlctr2_carry__2_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_5 ),
        .O(\i_sync_c[1]_i_346_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_347 
       (.I0(\I_0/hlctr2_carry__1_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_7 ),
        .O(\i_sync_c[1]_i_347_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_348 
       (.I0(\I_0/hlctr2_carry__1_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_5 ),
        .O(\i_sync_c[1]_i_348_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_349 
       (.I0(\I_0/hlctr2_carry__0_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_7 ),
        .O(\i_sync_c[1]_i_349_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_35 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_350 
       (.I0(\I_0/hlctr2_carry__2_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__2_n_6 ),
        .O(\i_sync_c[1]_i_350_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_351 
       (.I0(\I_0/hlctr2_carry__2_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_4 ),
        .O(\i_sync_c[1]_i_351_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_352 
       (.I0(\I_0/hlctr2_carry__1_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__1_n_6 ),
        .O(\i_sync_c[1]_i_352_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_353 
       (.I0(\I_0/hlctr2_carry__1_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_4 ),
        .O(\i_sync_c[1]_i_353_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_354 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_354_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_355 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_355_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_356 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_356_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_357 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_357_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_358 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_358_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_359 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_359_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_360 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_360_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_361 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_361_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_362 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_362_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_363 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_363_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_364 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_364_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_365 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_365_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_366 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_6 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_366_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_367 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_367_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_368 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_368_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \i_sync_c[1]_i_369 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_369_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_37 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_370 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_370_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_371 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_371_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_372 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_372_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_373 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_373_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_374 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_374_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_375 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_375_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h51)) 
    \i_sync_c[1]_i_376 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_376_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_377 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_377_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_378 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_378_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \i_sync_c[1]_i_379 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_379_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_38 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_380 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_380_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_381 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_381_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_382 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_382_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \i_sync_c[1]_i_383 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_383_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_384 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(\i_sync_c[1]_i_384_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_385 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_385_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_386 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_386_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_387 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_387_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \i_sync_c[1]_i_388 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_388_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_389 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_389_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_39 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \i_sync_c[1]_i_390 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_390_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_391 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_391_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_392 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_392_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_393 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_393_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_394 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(\i_sync_c[1]_i_394_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \i_sync_c[1]_i_395 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_395_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_396 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_396_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF7)) 
    \i_sync_c[1]_i_397 
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_397_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_398 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_398_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_399 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_4 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_399_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \i_sync_c[1]_i_4 
       (.I0(\I_0/i_sync_c218_in ),
        .I1(\I_0/i_sync_c219_in ),
        .O(\i_sync_c[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_40 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \i_sync_c[1]_i_400 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_400_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_401 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_401_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \i_sync_c[1]_i_402 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_402_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_403 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_403_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_404 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_404_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_405 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_405_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_406 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_7 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_406_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_407 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_407_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_408 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_408_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_409 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_409_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_41 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_410 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_410_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_411 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_411_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_412 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_4 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_412_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \i_sync_c[1]_i_413 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_413_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_414 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_414_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_415 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_415_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \i_sync_c[1]_i_416 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_416_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_417 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_417_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i_sync_c[1]_i_418 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_418_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_419 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_419_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_420 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_420_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_421 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_5 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_421_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \i_sync_c[1]_i_422 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_422_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_423 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_423_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_424 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_424_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_425 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_7 ),
        .I2(\I_0/hlctr_reg_n_0_ ),
        .O(\i_sync_c[1]_i_425_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_426 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_426_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_427 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_427_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_428 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_6 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_428_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h08)) 
    \i_sync_c[1]_i_429 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_429_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_43 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_430 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_430_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \i_sync_c[1]_i_431 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_431_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_432 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_432_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_433 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_433_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_434 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_434_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_435 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_435_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_436 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_6 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_436_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_437 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_437_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_438 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_438_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_439 
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_439_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_44 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_440 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_440_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_441 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__0_n_6 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_441_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \i_sync_c[1]_i_442 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_442_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_443 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_443_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \i_sync_c[1]_i_444 
       (.I0(\I_0/hlctr_reg_n_0_ ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_444_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_445 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_445_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_446 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_446_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_447 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_447_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_448 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry_n_6 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_448_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_449 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_449_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_45 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_450 
       (.I0(\I_0/hlctr2_carry__0_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_5 ),
        .O(\i_sync_c[1]_i_450_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_451 
       (.I0(\I_0/hlctr2_carry_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_7 ),
        .O(\i_sync_c[1]_i_451_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_452 
       (.I0(\I_0/hlctr2_carry_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_5 ),
        .O(\i_sync_c[1]_i_452_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h51)) 
    \i_sync_c[1]_i_453 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr2_carry_n_7 ),
        .O(\i_sync_c[1]_i_453_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_454 
       (.I0(\I_0/hlctr2_carry__0_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__0_n_6 ),
        .O(\i_sync_c[1]_i_454_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_455 
       (.I0(\I_0/hlctr2_carry__0_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_4 ),
        .O(\i_sync_c[1]_i_455_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_456 
       (.I0(\I_0/hlctr2_carry_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry_n_6 ),
        .O(\i_sync_c[1]_i_456_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \i_sync_c[1]_i_457 
       (.I0(\I_0/hlctr2_carry_n_7 ),
        .I1(\I_0/hlctr_reg_n_0_ ),
        .I2(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_457_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_46 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_47 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_48 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_49 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \i_sync_c[1]_i_5 
       (.I0(\I_0/i_sync_c229_in ),
        .I1(\I_0/i_sync_c28_in ),
        .O(\i_sync_c[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_50 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_52 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_53 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_54 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_55 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_56 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_57 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_58 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_59 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_61 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_62 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_63 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_64 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_65 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_66 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_67 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_68 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_70 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_71 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_72 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_73 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_74 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_76 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_77 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_78 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_79 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_80 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_82 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_83 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_84 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_85 
       (.I0(\I_0/hlctr2_carry__4_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_7 ),
        .O(\i_sync_c[1]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_86 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_87 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_88 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_89 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i_sync_c[1]_i_91 
       (.I0(\I_0/hlctr2_carry__6_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .O(\i_sync_c[1]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \i_sync_c[1]_i_92 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_93 
       (.I0(\I_0/hlctr2_carry__6_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_4 ),
        .O(\i_sync_c[1]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_94 
       (.I0(\I_0/hlctr2_carry__5_n_5 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_6 ),
        .O(\i_sync_c[1]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    \i_sync_c[1]_i_95 
       (.I0(\I_0/hlctr2_carry__5_n_7 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__4_n_4 ),
        .O(\i_sync_c[1]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    \i_sync_c[1]_i_97 
       (.I0(\I_0/hlctr1_carry__1_n_1 ),
        .I1(\I_0/hlctr2_carry__6_n_6 ),
        .I2(\I_0/hlctr2_carry__6_n_5 ),
        .O(\i_sync_c[1]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_98 
       (.I0(\I_0/hlctr2_carry__5_n_4 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__6_n_7 ),
        .O(\i_sync_c[1]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \i_sync_c[1]_i_99 
       (.I0(\I_0/hlctr2_carry__5_n_6 ),
        .I1(\I_0/hlctr1_carry__1_n_1 ),
        .I2(\I_0/hlctr2_carry__5_n_5 ),
        .O(\i_sync_c[1]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_10 
       (.CI(\i_sync_c_reg[1]_i_51_n_0 ),
        .CO({\I_0/i_sync_c224_in ,\i_sync_c_reg[1]_i_10_n_1 ,\i_sync_c_reg[1]_i_10_n_2 ,\i_sync_c_reg[1]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_52_n_0 ,\i_sync_c[1]_i_53_n_0 ,\i_sync_c[1]_i_54_n_0 ,\i_sync_c[1]_i_55_n_0 }),
        .S({\i_sync_c[1]_i_56_n_0 ,\i_sync_c[1]_i_57_n_0 ,\i_sync_c[1]_i_58_n_0 ,\i_sync_c[1]_i_59_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_105 
       (.CI(\i_sync_c_reg[1]_i_214_n_0 ),
        .CO(i_sync_c_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_215_n_0 ,\i_sync_c[1]_i_216_n_0 ,\i_sync_c[1]_i_217_n_0 ,\i_sync_c[1]_i_218_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_11 
       (.CI(\i_sync_c_reg[1]_i_60_n_0 ),
        .CO({\I_0/i_sync_c213_in ,\i_sync_c_reg[1]_i_11_n_1 ,\i_sync_c_reg[1]_i_11_n_2 ,\i_sync_c_reg[1]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_61_n_0 ,\i_sync_c[1]_i_62_n_0 ,\i_sync_c[1]_i_63_n_0 ,\i_sync_c[1]_i_64_n_0 }),
        .S({\i_sync_c[1]_i_65_n_0 ,\i_sync_c[1]_i_66_n_0 ,\i_sync_c[1]_i_67_n_0 ,\i_sync_c[1]_i_68_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_111 
       (.CI(\i_sync_c_reg[1]_i_219_n_0 ),
        .CO({\i_sync_c_reg[1]_i_111_n_0 ,\i_sync_c_reg[1]_i_111_n_1 ,\i_sync_c_reg[1]_i_111_n_2 ,\i_sync_c_reg[1]_i_111_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_220_n_0 ,\i_sync_c[1]_i_221_n_0 ,\i_sync_c[1]_i_222_n_0 ,\i_sync_c[1]_i_223_n_0 }),
        .S({\i_sync_c[1]_i_224_n_0 ,\i_sync_c[1]_i_225_n_0 ,\i_sync_c[1]_i_226_n_0 ,\i_sync_c[1]_i_227_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_12 
       (.CI(\i_sync_c_reg[1]_i_69_n_0 ),
        .CO({\I_0/i_sync_c212_in ,\i_sync_c_reg[1]_i_12_n_1 ,\i_sync_c_reg[1]_i_12_n_2 ,\i_sync_c_reg[1]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_70_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_71_n_0 ,\i_sync_c[1]_i_72_n_0 ,\i_sync_c[1]_i_73_n_0 ,\i_sync_c[1]_i_74_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_120 
       (.CI(\i_sync_c_reg[1]_i_228_n_0 ),
        .CO({\i_sync_c_reg[1]_i_120_n_0 ,\i_sync_c_reg[1]_i_120_n_1 ,\i_sync_c_reg[1]_i_120_n_2 ,\i_sync_c_reg[1]_i_120_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_229_n_0 ,\i_sync_c[1]_i_230_n_0 ,\i_sync_c[1]_i_231_n_0 ,\i_sync_c[1]_i_232_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_126 
       (.CI(\i_sync_c_reg[1]_i_233_n_0 ),
        .CO({\i_sync_c_reg[1]_i_126_n_0 ,\i_sync_c_reg[1]_i_126_n_1 ,\i_sync_c_reg[1]_i_126_n_2 ,\i_sync_c_reg[1]_i_126_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_234_n_0 ,\i_sync_c[1]_i_235_n_0 ,\i_sync_c[1]_i_236_n_0 ,\i_sync_c[1]_i_237_n_0 }),
        .S({\i_sync_c[1]_i_238_n_0 ,\i_sync_c[1]_i_239_n_0 ,\i_sync_c[1]_i_240_n_0 ,\i_sync_c[1]_i_241_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_13 
       (.CI(\i_sync_c_reg[1]_i_75_n_0 ),
        .CO({\I_0/i_sync_c210_in ,\i_sync_c_reg[1]_i_13_n_1 ,\i_sync_c_reg[1]_i_13_n_2 ,\i_sync_c_reg[1]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_76_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_77_n_0 ,\i_sync_c[1]_i_78_n_0 ,\i_sync_c[1]_i_79_n_0 ,\i_sync_c[1]_i_80_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_135 
       (.CI(\i_sync_c_reg[1]_i_242_n_0 ),
        .CO({\i_sync_c_reg[1]_i_135_n_0 ,\i_sync_c_reg[1]_i_135_n_1 ,\i_sync_c_reg[1]_i_135_n_2 ,\i_sync_c_reg[1]_i_135_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_243_n_0 ,\i_sync_c[1]_i_244_n_0 ,\i_sync_c[1]_i_245_n_0 ,\i_sync_c[1]_i_246_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_14 
       (.CI(\i_sync_c_reg[1]_i_81_n_0 ),
        .CO({\I_0/i_sync_c211_in ,\i_sync_c_reg[1]_i_14_n_1 ,\i_sync_c_reg[1]_i_14_n_2 ,\i_sync_c_reg[1]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_82_n_0 ,\i_sync_c[1]_i_83_n_0 ,\i_sync_c[1]_i_84_n_0 ,\i_sync_c[1]_i_85_n_0 }),
        .S({\i_sync_c[1]_i_86_n_0 ,\i_sync_c[1]_i_87_n_0 ,\i_sync_c[1]_i_88_n_0 ,\i_sync_c[1]_i_89_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_140 
       (.CI(\i_sync_c_reg[1]_i_247_n_0 ),
        .CO({\i_sync_c_reg[1]_i_140_n_0 ,\i_sync_c_reg[1]_i_140_n_1 ,\i_sync_c_reg[1]_i_140_n_2 ,\i_sync_c_reg[1]_i_140_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_248_n_0 ,\i_sync_c[1]_i_249_n_0 ,\i_sync_c[1]_i_250_n_0 ,\i_sync_c[1]_i_251_n_0 }),
        .S({\i_sync_c[1]_i_252_n_0 ,\i_sync_c[1]_i_253_n_0 ,\i_sync_c[1]_i_254_n_0 ,\i_sync_c[1]_i_255_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_149 
       (.CI(\i_sync_c_reg[1]_i_256_n_0 ),
        .CO({\i_sync_c_reg[1]_i_149_n_0 ,\i_sync_c_reg[1]_i_149_n_1 ,\i_sync_c_reg[1]_i_149_n_2 ,\i_sync_c_reg[1]_i_149_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_257_n_0 }),
        .S({\i_sync_c[1]_i_258_n_0 ,\i_sync_c[1]_i_259_n_0 ,\i_sync_c[1]_i_260_n_0 ,\i_sync_c[1]_i_261_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_15 
       (.CI(\i_sync_c_reg[1]_i_90_n_0 ),
        .CO({\I_0/i_sync_c215_in ,\i_sync_c_reg[1]_i_15_n_1 ,\i_sync_c_reg[1]_i_15_n_2 ,\i_sync_c_reg[1]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_91_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_92_n_0 ,\i_sync_c[1]_i_93_n_0 ,\i_sync_c[1]_i_94_n_0 ,\i_sync_c[1]_i_95_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_154 
       (.CI(\i_sync_c_reg[1]_i_262_n_0 ),
        .CO({\i_sync_c_reg[1]_i_154_n_0 ,\i_sync_c_reg[1]_i_154_n_1 ,\i_sync_c_reg[1]_i_154_n_2 ,\i_sync_c_reg[1]_i_154_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_263_n_0 ,\i_sync_c[1]_i_264_n_0 ,\i_sync_c[1]_i_265_n_0 ,\i_sync_c[1]_i_266_n_0 }),
        .S({\i_sync_c[1]_i_267_n_0 ,\i_sync_c[1]_i_268_n_0 ,\i_sync_c[1]_i_269_n_0 ,\i_sync_c[1]_i_270_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_16 
       (.CI(\i_sync_c_reg[1]_i_96_n_0 ),
        .CO({\I_0/i_sync_c216_in ,\i_sync_c_reg[1]_i_16_n_1 ,\i_sync_c_reg[1]_i_16_n_2 ,\i_sync_c_reg[1]_i_16_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_97_n_0 ,\i_sync_c[1]_i_98_n_0 ,\i_sync_c[1]_i_99_n_0 ,\i_sync_c[1]_i_100_n_0 }),
        .S({\i_sync_c[1]_i_101_n_0 ,\i_sync_c[1]_i_102_n_0 ,\i_sync_c[1]_i_103_n_0 ,\i_sync_c[1]_i_104_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_163 
       (.CI(\i_sync_c_reg[1]_i_271_n_0 ),
        .CO({\i_sync_c_reg[1]_i_163_n_0 ,\i_sync_c_reg[1]_i_163_n_1 ,\i_sync_c_reg[1]_i_163_n_2 ,\i_sync_c_reg[1]_i_163_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_272_n_0 ,\i_sync_c[1]_i_273_n_0 ,\i_sync_c[1]_i_274_n_0 ,\i_sync_c[1]_i_275_n_0 }),
        .S({\i_sync_c[1]_i_276_n_0 ,\i_sync_c[1]_i_277_n_0 ,\i_sync_c[1]_i_278_n_0 ,\i_sync_c[1]_i_279_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_17 
       (.CI(i_sync_c_reg[3]),
        .CO({\I_0/i_sync_c218_in ,\i_sync_c_reg[1]_i_17_n_1 ,\i_sync_c_reg[1]_i_17_n_2 ,\i_sync_c_reg[1]_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_106_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_107_n_0 ,\i_sync_c[1]_i_108_n_0 ,\i_sync_c[1]_i_109_n_0 ,\i_sync_c[1]_i_110_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_172 
       (.CI(\i_sync_c_reg[1]_i_280_n_0 ),
        .CO({\i_sync_c_reg[1]_i_172_n_0 ,\i_sync_c_reg[1]_i_172_n_1 ,\i_sync_c_reg[1]_i_172_n_2 ,\i_sync_c_reg[1]_i_172_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_281_n_0 ,\i_sync_c[1]_i_282_n_0 ,\i_sync_c[1]_i_283_n_0 ,\i_sync_c[1]_i_284_n_0 }),
        .S({\i_sync_c[1]_i_285_n_0 ,\i_sync_c[1]_i_286_n_0 ,\i_sync_c[1]_i_287_n_0 ,\i_sync_c[1]_i_288_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_18 
       (.CI(\i_sync_c_reg[1]_i_111_n_0 ),
        .CO({\I_0/i_sync_c219_in ,\i_sync_c_reg[1]_i_18_n_1 ,\i_sync_c_reg[1]_i_18_n_2 ,\i_sync_c_reg[1]_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_112_n_0 ,\i_sync_c[1]_i_113_n_0 ,\i_sync_c[1]_i_114_n_0 ,\i_sync_c[1]_i_115_n_0 }),
        .S({\i_sync_c[1]_i_116_n_0 ,\i_sync_c[1]_i_117_n_0 ,\i_sync_c[1]_i_118_n_0 ,\i_sync_c[1]_i_119_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_181 
       (.CI(\i_sync_c_reg[1]_i_289_n_0 ),
        .CO({\i_sync_c_reg[1]_i_181_n_0 ,\i_sync_c_reg[1]_i_181_n_1 ,\i_sync_c_reg[1]_i_181_n_2 ,\i_sync_c_reg[1]_i_181_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_290_n_0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_291_n_0 ,\i_sync_c[1]_i_292_n_0 ,\i_sync_c[1]_i_293_n_0 ,\i_sync_c[1]_i_294_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_186 
       (.CI(\i_sync_c_reg[1]_i_295_n_0 ),
        .CO({\i_sync_c_reg[1]_i_186_n_0 ,\i_sync_c_reg[1]_i_186_n_1 ,\i_sync_c_reg[1]_i_186_n_2 ,\i_sync_c_reg[1]_i_186_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_296_n_0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_297_n_0 ,\i_sync_c[1]_i_298_n_0 ,\i_sync_c[1]_i_299_n_0 ,\i_sync_c[1]_i_300_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_19 
       (.CI(\i_sync_c_reg[1]_i_120_n_0 ),
        .CO({\I_0/i_sync_c229_in ,\i_sync_c_reg[1]_i_19_n_1 ,\i_sync_c_reg[1]_i_19_n_2 ,\i_sync_c_reg[1]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_121_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_122_n_0 ,\i_sync_c[1]_i_123_n_0 ,\i_sync_c[1]_i_124_n_0 ,\i_sync_c[1]_i_125_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_191 
       (.CI(\i_sync_c_reg[1]_i_301_n_0 ),
        .CO({\i_sync_c_reg[1]_i_191_n_0 ,\i_sync_c_reg[1]_i_191_n_1 ,\i_sync_c_reg[1]_i_191_n_2 ,\i_sync_c_reg[1]_i_191_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_302_n_0 ,\i_sync_c[1]_i_303_n_0 ,\i_sync_c[1]_i_304_n_0 ,\i_sync_c[1]_i_305_n_0 }),
        .S({\i_sync_c[1]_i_306_n_0 ,\i_sync_c[1]_i_307_n_0 ,\i_sync_c[1]_i_308_n_0 ,\i_sync_c[1]_i_309_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_20 
       (.CI(\i_sync_c_reg[1]_i_126_n_0 ),
        .CO({\I_0/i_sync_c28_in ,\i_sync_c_reg[1]_i_20_n_1 ,\i_sync_c_reg[1]_i_20_n_2 ,\i_sync_c_reg[1]_i_20_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_127_n_0 ,\i_sync_c[1]_i_128_n_0 ,\i_sync_c[1]_i_129_n_0 ,\i_sync_c[1]_i_130_n_0 }),
        .S({\i_sync_c[1]_i_131_n_0 ,\i_sync_c[1]_i_132_n_0 ,\i_sync_c[1]_i_133_n_0 ,\i_sync_c[1]_i_134_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_200 
       (.CI(\i_sync_c_reg[1]_i_310_n_0 ),
        .CO({\i_sync_c_reg[1]_i_200_n_0 ,\i_sync_c_reg[1]_i_200_n_1 ,\i_sync_c_reg[1]_i_200_n_2 ,\i_sync_c_reg[1]_i_200_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_311_n_0 }),
        .S({\i_sync_c[1]_i_312_n_0 ,\i_sync_c[1]_i_313_n_0 ,\i_sync_c[1]_i_314_n_0 ,\i_sync_c[1]_i_315_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_205 
       (.CI(\i_sync_c_reg[1]_i_316_n_0 ),
        .CO({\i_sync_c_reg[1]_i_205_n_0 ,\i_sync_c_reg[1]_i_205_n_1 ,\i_sync_c_reg[1]_i_205_n_2 ,\i_sync_c_reg[1]_i_205_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_317_n_0 ,\i_sync_c[1]_i_318_n_0 ,\i_sync_c[1]_i_319_n_0 ,\i_sync_c[1]_i_320_n_0 }),
        .S({\i_sync_c[1]_i_321_n_0 ,\i_sync_c[1]_i_322_n_0 ,\i_sync_c[1]_i_323_n_0 ,\i_sync_c[1]_i_324_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_21 
       (.CI(\i_sync_c_reg[1]_i_135_n_0 ),
        .CO({\i_sync_c_reg[1]_i_21_n_0 ,\i_sync_c_reg[1]_i_21_n_1 ,\i_sync_c_reg[1]_i_21_n_2 ,\i_sync_c_reg[1]_i_21_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_136_n_0 ,\i_sync_c[1]_i_137_n_0 ,\i_sync_c[1]_i_138_n_0 ,\i_sync_c[1]_i_139_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_214 
       (.CI(\i_sync_c_reg[1]_i_325_n_0 ),
        .CO({\i_sync_c_reg[1]_i_214_n_0 ,\i_sync_c_reg[1]_i_214_n_1 ,\i_sync_c_reg[1]_i_214_n_2 ,\i_sync_c_reg[1]_i_214_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_326_n_0 }),
        .S({\i_sync_c[1]_i_327_n_0 ,\i_sync_c[1]_i_328_n_0 ,\i_sync_c[1]_i_329_n_0 ,\i_sync_c[1]_i_330_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_219 
       (.CI(\i_sync_c_reg[1]_i_331_n_0 ),
        .CO({\i_sync_c_reg[1]_i_219_n_0 ,\i_sync_c_reg[1]_i_219_n_1 ,\i_sync_c_reg[1]_i_219_n_2 ,\i_sync_c_reg[1]_i_219_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_332_n_0 ,\i_sync_c[1]_i_333_n_0 ,\i_sync_c[1]_i_334_n_0 ,\i_sync_c[1]_i_335_n_0 }),
        .S({\i_sync_c[1]_i_336_n_0 ,\i_sync_c[1]_i_337_n_0 ,\i_sync_c[1]_i_338_n_0 ,\i_sync_c[1]_i_339_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_228 
       (.CI(\i_sync_c_reg[1]_i_340_n_0 ),
        .CO({\i_sync_c_reg[1]_i_228_n_0 ,\i_sync_c_reg[1]_i_228_n_1 ,\i_sync_c_reg[1]_i_228_n_2 ,\i_sync_c_reg[1]_i_228_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_341_n_0 ,\i_sync_c[1]_i_342_n_0 ,\i_sync_c[1]_i_343_n_0 ,\i_sync_c[1]_i_344_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_233 
       (.CI(\i_sync_c_reg[1]_i_345_n_0 ),
        .CO({\i_sync_c_reg[1]_i_233_n_0 ,\i_sync_c_reg[1]_i_233_n_1 ,\i_sync_c_reg[1]_i_233_n_2 ,\i_sync_c_reg[1]_i_233_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_346_n_0 ,\i_sync_c[1]_i_347_n_0 ,\i_sync_c[1]_i_348_n_0 ,\i_sync_c[1]_i_349_n_0 }),
        .S({\i_sync_c[1]_i_350_n_0 ,\i_sync_c[1]_i_351_n_0 ,\i_sync_c[1]_i_352_n_0 ,\i_sync_c[1]_i_353_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_242 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_242_n_0 ,\i_sync_c_reg[1]_i_242_n_1 ,\i_sync_c_reg[1]_i_242_n_2 ,\i_sync_c_reg[1]_i_242_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_354_n_0 ,\i_sync_c[1]_i_355_n_0 }),
        .S({\i_sync_c[1]_i_356_n_0 ,\i_sync_c[1]_i_357_n_0 ,\i_sync_c[1]_i_358_n_0 ,\i_sync_c[1]_i_359_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_247 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_247_n_0 ,\i_sync_c_reg[1]_i_247_n_1 ,\i_sync_c_reg[1]_i_247_n_2 ,\i_sync_c_reg[1]_i_247_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_360_n_0 ,\i_sync_c[1]_i_361_n_0 ,\i_sync_c[1]_i_362_n_0 ,\i_sync_c[1]_i_363_n_0 }),
        .S({\i_sync_c[1]_i_364_n_0 ,\i_sync_c[1]_i_365_n_0 ,\i_sync_c[1]_i_366_n_0 ,\i_sync_c[1]_i_367_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_256 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_256_n_0 ,\i_sync_c_reg[1]_i_256_n_1 ,\i_sync_c_reg[1]_i_256_n_2 ,\i_sync_c_reg[1]_i_256_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_368_n_0 ,\i_sync_c[1]_i_369_n_0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_370_n_0 ,\i_sync_c[1]_i_371_n_0 ,\i_sync_c[1]_i_372_n_0 ,\i_sync_c[1]_i_373_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_262 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_262_n_0 ,\i_sync_c_reg[1]_i_262_n_1 ,\i_sync_c_reg[1]_i_262_n_2 ,\i_sync_c_reg[1]_i_262_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_374_n_0 ,\i_sync_c[1]_i_375_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_376_n_0 }),
        .S({\i_sync_c[1]_i_377_n_0 ,\i_sync_c[1]_i_378_n_0 ,\i_sync_c[1]_i_379_n_0 ,\i_sync_c[1]_i_380_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_27 
       (.CI(\i_sync_c_reg[1]_i_140_n_0 ),
        .CO({\i_sync_c_reg[1]_i_27_n_0 ,\i_sync_c_reg[1]_i_27_n_1 ,\i_sync_c_reg[1]_i_27_n_2 ,\i_sync_c_reg[1]_i_27_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_141_n_0 ,\i_sync_c[1]_i_142_n_0 ,\i_sync_c[1]_i_143_n_0 ,\i_sync_c[1]_i_144_n_0 }),
        .S({\i_sync_c[1]_i_145_n_0 ,\i_sync_c[1]_i_146_n_0 ,\i_sync_c[1]_i_147_n_0 ,\i_sync_c[1]_i_148_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_271 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_271_n_0 ,\i_sync_c_reg[1]_i_271_n_1 ,\i_sync_c_reg[1]_i_271_n_2 ,\i_sync_c_reg[1]_i_271_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_381_n_0 ,\i_sync_c[1]_i_382_n_0 ,\i_sync_c[1]_i_383_n_0 ,\i_sync_c[1]_i_384_n_0 }),
        .S({\i_sync_c[1]_i_385_n_0 ,\i_sync_c[1]_i_386_n_0 ,\i_sync_c[1]_i_387_n_0 ,\i_sync_c[1]_i_388_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_280 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_280_n_0 ,\i_sync_c_reg[1]_i_280_n_1 ,\i_sync_c_reg[1]_i_280_n_2 ,\i_sync_c_reg[1]_i_280_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_389_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_390_n_0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_391_n_0 ,\i_sync_c[1]_i_392_n_0 ,\i_sync_c[1]_i_393_n_0 ,\i_sync_c[1]_i_394_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_289 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_289_n_0 ,\i_sync_c_reg[1]_i_289_n_1 ,\i_sync_c_reg[1]_i_289_n_2 ,\i_sync_c_reg[1]_i_289_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_395_n_0 ,\i_sync_c[1]_i_396_n_0 ,\i_sync_c[1]_i_397_n_0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_398_n_0 ,\i_sync_c[1]_i_399_n_0 ,\i_sync_c[1]_i_400_n_0 ,\i_sync_c[1]_i_401_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_295 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_295_n_0 ,\i_sync_c_reg[1]_i_295_n_1 ,\i_sync_c_reg[1]_i_295_n_2 ,\i_sync_c_reg[1]_i_295_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_402_n_0 ,\i_sync_c[1]_i_403_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_404_n_0 }),
        .S({\i_sync_c[1]_i_405_n_0 ,\i_sync_c[1]_i_406_n_0 ,\i_sync_c[1]_i_407_n_0 ,\i_sync_c[1]_i_408_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_301 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_301_n_0 ,\i_sync_c_reg[1]_i_301_n_1 ,\i_sync_c_reg[1]_i_301_n_2 ,\i_sync_c_reg[1]_i_301_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\i_sync_c[1]_i_409_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_410_n_0 }),
        .S({\i_sync_c[1]_i_411_n_0 ,\i_sync_c[1]_i_412_n_0 ,\i_sync_c[1]_i_413_n_0 ,\i_sync_c[1]_i_414_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_310 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_310_n_0 ,\i_sync_c_reg[1]_i_310_n_1 ,\i_sync_c_reg[1]_i_310_n_2 ,\i_sync_c_reg[1]_i_310_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_415_n_0 ,\i_sync_c[1]_i_416_n_0 ,\i_sync_c[1]_i_417_n_0 ,\i_sync_c[1]_i_418_n_0 }),
        .S({\i_sync_c[1]_i_419_n_0 ,\i_sync_c[1]_i_420_n_0 ,\i_sync_c[1]_i_421_n_0 ,\i_sync_c[1]_i_422_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_316 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_316_n_0 ,\i_sync_c_reg[1]_i_316_n_1 ,\i_sync_c_reg[1]_i_316_n_2 ,\i_sync_c_reg[1]_i_316_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_423_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_424_n_0 ,\i_sync_c[1]_i_425_n_0 }),
        .S({\i_sync_c[1]_i_426_n_0 ,\i_sync_c[1]_i_427_n_0 ,\i_sync_c[1]_i_428_n_0 ,\i_sync_c[1]_i_429_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_325 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_325_n_0 ,\i_sync_c_reg[1]_i_325_n_1 ,\i_sync_c_reg[1]_i_325_n_2 ,\i_sync_c_reg[1]_i_325_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_430_n_0 ,\i_sync_c[1]_i_431_n_0 ,\i_sync_c[1]_i_432_n_0 ,\i_sync_c[1]_i_433_n_0 }),
        .S({\i_sync_c[1]_i_434_n_0 ,\i_sync_c[1]_i_435_n_0 ,\i_sync_c[1]_i_436_n_0 ,\i_sync_c[1]_i_437_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_331 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_331_n_0 ,\i_sync_c_reg[1]_i_331_n_1 ,\i_sync_c_reg[1]_i_331_n_2 ,\i_sync_c_reg[1]_i_331_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_438_n_0 ,\<const0>__0__0 ,\i_sync_c[1]_i_439_n_0 ,\i_sync_c[1]_i_440_n_0 }),
        .S({\i_sync_c[1]_i_441_n_0 ,\i_sync_c[1]_i_442_n_0 ,\i_sync_c[1]_i_443_n_0 ,\i_sync_c[1]_i_444_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_340 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_340_n_0 ,\i_sync_c_reg[1]_i_340_n_1 ,\i_sync_c_reg[1]_i_340_n_2 ,\i_sync_c_reg[1]_i_340_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\i_sync_c[1]_i_445_n_0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_446_n_0 ,\i_sync_c[1]_i_447_n_0 ,\i_sync_c[1]_i_448_n_0 ,\i_sync_c[1]_i_449_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_345 
       (.CI(\<const0>__0__0 ),
        .CO({\i_sync_c_reg[1]_i_345_n_0 ,\i_sync_c_reg[1]_i_345_n_1 ,\i_sync_c_reg[1]_i_345_n_2 ,\i_sync_c_reg[1]_i_345_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\i_sync_c[1]_i_450_n_0 ,\i_sync_c[1]_i_451_n_0 ,\i_sync_c[1]_i_452_n_0 ,\i_sync_c[1]_i_453_n_0 }),
        .S({\i_sync_c[1]_i_454_n_0 ,\i_sync_c[1]_i_455_n_0 ,\i_sync_c[1]_i_456_n_0 ,\i_sync_c[1]_i_457_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_36 
       (.CI(\i_sync_c_reg[1]_i_149_n_0 ),
        .CO({\i_sync_c_reg[1]_i_36_n_0 ,\i_sync_c_reg[1]_i_36_n_1 ,\i_sync_c_reg[1]_i_36_n_2 ,\i_sync_c_reg[1]_i_36_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_150_n_0 ,\i_sync_c[1]_i_151_n_0 ,\i_sync_c[1]_i_152_n_0 ,\i_sync_c[1]_i_153_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_42 
       (.CI(\i_sync_c_reg[1]_i_154_n_0 ),
        .CO({\i_sync_c_reg[1]_i_42_n_0 ,\i_sync_c_reg[1]_i_42_n_1 ,\i_sync_c_reg[1]_i_42_n_2 ,\i_sync_c_reg[1]_i_42_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_155_n_0 ,\i_sync_c[1]_i_156_n_0 ,\i_sync_c[1]_i_157_n_0 ,\i_sync_c[1]_i_158_n_0 }),
        .S({\i_sync_c[1]_i_159_n_0 ,\i_sync_c[1]_i_160_n_0 ,\i_sync_c[1]_i_161_n_0 ,\i_sync_c[1]_i_162_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_51 
       (.CI(\i_sync_c_reg[1]_i_163_n_0 ),
        .CO({\i_sync_c_reg[1]_i_51_n_0 ,\i_sync_c_reg[1]_i_51_n_1 ,\i_sync_c_reg[1]_i_51_n_2 ,\i_sync_c_reg[1]_i_51_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_164_n_0 ,\i_sync_c[1]_i_165_n_0 ,\i_sync_c[1]_i_166_n_0 ,\i_sync_c[1]_i_167_n_0 }),
        .S({\i_sync_c[1]_i_168_n_0 ,\i_sync_c[1]_i_169_n_0 ,\i_sync_c[1]_i_170_n_0 ,\i_sync_c[1]_i_171_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_6 
       (.CI(\i_sync_c_reg[1]_i_21_n_0 ),
        .CO({\I_0/i_sync_c226_in ,\i_sync_c_reg[1]_i_6_n_1 ,\i_sync_c_reg[1]_i_6_n_2 ,\i_sync_c_reg[1]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_22_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_23_n_0 ,\i_sync_c[1]_i_24_n_0 ,\i_sync_c[1]_i_25_n_0 ,\i_sync_c[1]_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_60 
       (.CI(\i_sync_c_reg[1]_i_172_n_0 ),
        .CO({\i_sync_c_reg[1]_i_60_n_0 ,\i_sync_c_reg[1]_i_60_n_1 ,\i_sync_c_reg[1]_i_60_n_2 ,\i_sync_c_reg[1]_i_60_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_173_n_0 ,\i_sync_c[1]_i_174_n_0 ,\i_sync_c[1]_i_175_n_0 ,\i_sync_c[1]_i_176_n_0 }),
        .S({\i_sync_c[1]_i_177_n_0 ,\i_sync_c[1]_i_178_n_0 ,\i_sync_c[1]_i_179_n_0 ,\i_sync_c[1]_i_180_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_69 
       (.CI(\i_sync_c_reg[1]_i_181_n_0 ),
        .CO({\i_sync_c_reg[1]_i_69_n_0 ,\i_sync_c_reg[1]_i_69_n_1 ,\i_sync_c_reg[1]_i_69_n_2 ,\i_sync_c_reg[1]_i_69_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_182_n_0 ,\i_sync_c[1]_i_183_n_0 ,\i_sync_c[1]_i_184_n_0 ,\i_sync_c[1]_i_185_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_7 
       (.CI(\i_sync_c_reg[1]_i_27_n_0 ),
        .CO({\I_0/i_sync_c227_in ,\i_sync_c_reg[1]_i_7_n_1 ,\i_sync_c_reg[1]_i_7_n_2 ,\i_sync_c_reg[1]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_28_n_0 ,\i_sync_c[1]_i_29_n_0 ,\i_sync_c[1]_i_30_n_0 ,\i_sync_c[1]_i_31_n_0 }),
        .S({\i_sync_c[1]_i_32_n_0 ,\i_sync_c[1]_i_33_n_0 ,\i_sync_c[1]_i_34_n_0 ,\i_sync_c[1]_i_35_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_75 
       (.CI(\i_sync_c_reg[1]_i_186_n_0 ),
        .CO({\i_sync_c_reg[1]_i_75_n_0 ,\i_sync_c_reg[1]_i_75_n_1 ,\i_sync_c_reg[1]_i_75_n_2 ,\i_sync_c_reg[1]_i_75_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_187_n_0 ,\i_sync_c[1]_i_188_n_0 ,\i_sync_c[1]_i_189_n_0 ,\i_sync_c[1]_i_190_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_8 
       (.CI(\i_sync_c_reg[1]_i_36_n_0 ),
        .CO({\I_0/i_sync_c221_in ,\i_sync_c_reg[1]_i_8_n_1 ,\i_sync_c_reg[1]_i_8_n_2 ,\i_sync_c_reg[1]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_37_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_38_n_0 ,\i_sync_c[1]_i_39_n_0 ,\i_sync_c[1]_i_40_n_0 ,\i_sync_c[1]_i_41_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_81 
       (.CI(\i_sync_c_reg[1]_i_191_n_0 ),
        .CO({\i_sync_c_reg[1]_i_81_n_0 ,\i_sync_c_reg[1]_i_81_n_1 ,\i_sync_c_reg[1]_i_81_n_2 ,\i_sync_c_reg[1]_i_81_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_192_n_0 ,\i_sync_c[1]_i_193_n_0 ,\i_sync_c[1]_i_194_n_0 ,\i_sync_c[1]_i_195_n_0 }),
        .S({\i_sync_c[1]_i_196_n_0 ,\i_sync_c[1]_i_197_n_0 ,\i_sync_c[1]_i_198_n_0 ,\i_sync_c[1]_i_199_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_9 
       (.CI(\i_sync_c_reg[1]_i_42_n_0 ),
        .CO({\I_0/i_sync_c2 ,\i_sync_c_reg[1]_i_9_n_1 ,\i_sync_c_reg[1]_i_9_n_2 ,\i_sync_c_reg[1]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_43_n_0 ,\i_sync_c[1]_i_44_n_0 ,\i_sync_c[1]_i_45_n_0 ,\i_sync_c[1]_i_46_n_0 }),
        .S({\i_sync_c[1]_i_47_n_0 ,\i_sync_c[1]_i_48_n_0 ,\i_sync_c[1]_i_49_n_0 ,\i_sync_c[1]_i_50_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_90 
       (.CI(\i_sync_c_reg[1]_i_200_n_0 ),
        .CO({\i_sync_c_reg[1]_i_90_n_0 ,\i_sync_c_reg[1]_i_90_n_1 ,\i_sync_c_reg[1]_i_90_n_2 ,\i_sync_c_reg[1]_i_90_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\i_sync_c[1]_i_201_n_0 ,\i_sync_c[1]_i_202_n_0 ,\i_sync_c[1]_i_203_n_0 ,\i_sync_c[1]_i_204_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \i_sync_c_reg[1]_i_96 
       (.CI(\i_sync_c_reg[1]_i_205_n_0 ),
        .CO({\i_sync_c_reg[1]_i_96_n_0 ,\i_sync_c_reg[1]_i_96_n_1 ,\i_sync_c_reg[1]_i_96_n_2 ,\i_sync_c_reg[1]_i_96_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\i_sync_c[1]_i_206_n_0 ,\i_sync_c[1]_i_207_n_0 ,\i_sync_c[1]_i_208_n_0 ,\i_sync_c[1]_i_209_n_0 }),
        .S({\i_sync_c[1]_i_210_n_0 ,\i_sync_c[1]_i_211_n_0 ,\i_sync_c[1]_i_212_n_0 ,\i_sync_c[1]_i_213_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_carry__0_i_1
       (.I0(in_r[3]),
        .I1(plusOp18[8]),
        .O(minusOp_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_carry__0_i_2
       (.I0(in_r[2]),
        .I1(plusOp18[7]),
        .O(minusOp_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_carry__0_i_3
       (.I0(in_r[1]),
        .I1(plusOp18[6]),
        .O(minusOp_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_carry__0_i_4
       (.I0(in_r[0]),
        .I1(plusOp18[5]),
        .O(minusOp_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_carry__1_i_2
       (.I0(in_r[4]),
        .I1(plusOp18[9]),
        .O(minusOp_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_1
       (.I0(in_b[3]),
        .I1(plusOp18[8]),
        .O(minusOp_inferred__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_2
       (.I0(in_b[2]),
        .I1(plusOp18[7]),
        .O(minusOp_inferred__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_3
       (.I0(in_b[1]),
        .I1(plusOp18[6]),
        .O(minusOp_inferred__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__0_i_4
       (.I0(in_b[0]),
        .I1(plusOp18[5]),
        .O(minusOp_inferred__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    minusOp_inferred__0_carry__1_i_2
       (.I0(in_b[4]),
        .I1(plusOp18[9]),
        .O(minusOp_inferred__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(1),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    modu_reg
       (.A({\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[15] ,\I_1/data_reg_n_0_[14] ,\I_1/data_reg_n_0_[13] ,\I_1/data_reg_n_0_[12] ,\I_1/data_reg_n_0_[11] ,\I_1/data_reg_n_0_[10] ,\I_1/data_reg_n_0_[9] ,\I_1/data_reg_n_0_[8] ,\I_1/data_reg_n_0_[7] ,\I_1/data_reg_n_0_[6] ,\I_1/data_reg_n_0_[5] ,\I_1/data_reg_n_0_[4] ,\I_1/data_reg_n_0_[3] ,\I_1/data_reg_n_0_[2] ,\I_1/data_reg_n_0_[1] ,\I_1/data_reg_n_0_ }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[11] ,\I_4/output_reg_n_0_[10] ,\I_4/output_reg_n_0_[9] ,\I_4/output_reg_n_0_[8] ,\I_4/output_reg_n_0_[7] ,\I_4/output_reg_n_0_[6] ,\I_4/output_reg_n_0_[5] ,\I_4/output_reg_n_0_[4] ,\I_4/output_reg_n_0_[3] ,\I_4/output_reg_n_0_[2] ,\I_4/output_reg_n_0_[1] ,\I_4/output_reg_n_0_ }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(reset),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({modu_reg_n_58,modu_reg_n_59,modu_reg_n_60,modu_reg_n_61,modu_reg_n_62,modu_reg_n_63,modu_reg_n_64,modu_reg_n_65,modu_reg_n_66,modu_reg_n_67,modu_reg_n_68,modu_reg_n_69,modu_reg_n_70,modu_reg_n_71,modu_reg_n_72,modu_reg_n_73,modu_reg_n_74,modu_reg_n_75,modu_reg_n_76,modu_reg_n_77,modu_reg_n_78,modu_reg_n_79,modu_reg_n_80,modu_reg_n_81,modu_reg_n_82,modu_reg_n_83,modu_reg_n_84,modu_reg_n_85,modu_reg_n_86,modu_reg_n_87,modu_reg_n_88,modu_reg_n_89,modu_reg_n_90,modu_reg_n_91,modu_reg_n_92,modu_reg_n_93,modu_reg_n_94,modu_reg_n_95,modu_reg_n_96,modu_reg_n_97,modu_reg_n_98,modu_reg_n_99,modu_reg_n_100,modu_reg_n_101,modu_reg_n_102,modu_reg_n_103,modu_reg_n_104,modu_reg_n_105}),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(1),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    modus_reg
       (.A({modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_79,modu_reg_n_80,modu_reg_n_81,modu_reg_n_82,modu_reg_n_83,modu_reg_n_84,modu_reg_n_85,modu_reg_n_86,modu_reg_n_87,modu_reg_n_88,modu_reg_n_89,modu_reg_n_90}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(reset),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({modus_reg_n_58,modus_reg_n_59,modus_reg_n_60,modus_reg_n_61,modus_reg_n_62,modus_reg_n_63,modus_reg_n_64,modus_reg_n_65,modus_reg_n_66,modus_reg_n_67,modus_reg_n_68,modus_reg_n_69,modus_reg_n_70,modus_reg_n_71,modus_reg_n_72,modus_reg_n_73,modus_reg_n_74,modus_reg_n_75,modus_reg_n_76,modus_reg_n_77,modus_reg_n_78,modus_reg_n_79,L,modus_reg_n_96,modus_reg_n_97,modus_reg_n_98,modus_reg_n_99,modus_reg_n_100,modus_reg_n_101,modus_reg_n_102,modus_reg_n_103,modus_reg_n_104,modus_reg_n_105}),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(1),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    modv_reg
       (.A({modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_1_n_0,modv_reg_i_2_n_0,modv_reg_i_3_n_0,modv_reg_i_4_n_0,modv_reg_i_5_n_0,modv_reg_i_6_n_0,modv_reg_i_7_n_0,modv_reg_i_8_n_0,modv_reg_i_9_n_0,modv_reg_i_10_n_0,modv_reg_i_11_n_0,modv_reg_i_12_n_0,modv_reg_i_13_n_0,modv_reg_i_14_n_0,modv_reg_i_15_n_0,data[0]}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[11] ,\I_5/output_reg_n_0_[10] ,\I_5/output_reg_n_0_[9] ,\I_5/output_reg_n_0_[8] ,\I_5/output_reg_n_0_[7] ,\I_5/output_reg_n_0_[6] ,\I_5/output_reg_n_0_[5] ,\I_5/output_reg_n_0_[4] ,\I_5/output_reg_n_0_[3] ,\I_5/output_reg_n_0_[2] ,\I_5/output_reg_n_0_[1] ,\I_5/output_reg_n_0_ }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(reset),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({modv_reg_n_58,modv_reg_n_59,modv_reg_n_60,modv_reg_n_61,modv_reg_n_62,modv_reg_n_63,modv_reg_n_64,modv_reg_n_65,modv_reg_n_66,modv_reg_n_67,modv_reg_n_68,modv_reg_n_69,modv_reg_n_70,modv_reg_n_71,modv_reg_n_72,modv_reg_n_73,modv_reg_n_74,modv_reg_n_75,modv_reg_n_76,modv_reg_n_77,modv_reg_n_78,A,modv_reg_n_91,modv_reg_n_92,modv_reg_n_93,modv_reg_n_94,modv_reg_n_95,modv_reg_n_96,modv_reg_n_97,modv_reg_n_98,modv_reg_n_99,modv_reg_n_100,modv_reg_n_101,modv_reg_n_102,modv_reg_n_103,modv_reg_n_104,modv_reg_n_105}),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_1
       (.I0(psin0[15]),
        .I1(phase),
        .I2(data[15]),
        .O(modv_reg_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_10
       (.I0(psin0[6]),
        .I1(phase),
        .I2(data[6]),
        .O(modv_reg_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_11
       (.I0(psin0[5]),
        .I1(phase),
        .I2(data[5]),
        .O(modv_reg_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_12
       (.I0(psin0[4]),
        .I1(phase),
        .I2(data[4]),
        .O(modv_reg_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_13
       (.I0(psin0[3]),
        .I1(phase),
        .I2(data[3]),
        .O(modv_reg_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_14
       (.I0(psin0[2]),
        .I1(phase),
        .I2(data[2]),
        .O(modv_reg_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_15
       (.I0(psin0[1]),
        .I1(phase),
        .I2(data[1]),
        .O(modv_reg_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 modv_reg_i_16
       (.CI(modv_reg_i_17_n_0),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({modv_reg_i_16_n_4,psin0[15:13]}),
        .S({\<const0>__0__0 ,modv_reg_i_20_n_0,modv_reg_i_21_n_0,modv_reg_i_22_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 modv_reg_i_17
       (.CI(modv_reg_i_18_n_0),
        .CO({modv_reg_i_17_n_0,modv_reg_i_17_n_1,modv_reg_i_17_n_2,modv_reg_i_17_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(psin0[12:9]),
        .S({modv_reg_i_23_n_0,modv_reg_i_24_n_0,modv_reg_i_25_n_0,modv_reg_i_26_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 modv_reg_i_18
       (.CI(modv_reg_i_19_n_0),
        .CO({modv_reg_i_18_n_0,modv_reg_i_18_n_1,modv_reg_i_18_n_2,modv_reg_i_18_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(psin0[8:5]),
        .S({modv_reg_i_27_n_0,modv_reg_i_28_n_0,modv_reg_i_29_n_0,modv_reg_i_30_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 modv_reg_i_19
       (.CI(\<const0>__0__0 ),
        .CO({modv_reg_i_19_n_0,modv_reg_i_19_n_1,modv_reg_i_19_n_2,modv_reg_i_19_n_3}),
        .CYINIT(modv_reg_i_31_n_0),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(psin0[4:1]),
        .S({modv_reg_i_32_n_0,modv_reg_i_33_n_0,modv_reg_i_34_n_0,modv_reg_i_35_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_2
       (.I0(psin0[14]),
        .I1(phase),
        .I2(data[14]),
        .O(modv_reg_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_20
       (.I0(data[15]),
        .O(modv_reg_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_21
       (.I0(data[14]),
        .O(modv_reg_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_22
       (.I0(data[13]),
        .O(modv_reg_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_23
       (.I0(data[12]),
        .O(modv_reg_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_24
       (.I0(data[11]),
        .O(modv_reg_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_25
       (.I0(data[10]),
        .O(modv_reg_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_26
       (.I0(data[9]),
        .O(modv_reg_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_27
       (.I0(data[8]),
        .O(modv_reg_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_28
       (.I0(data[7]),
        .O(modv_reg_i_28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_29
       (.I0(data[6]),
        .O(modv_reg_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_3
       (.I0(psin0[13]),
        .I1(phase),
        .I2(data[13]),
        .O(modv_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_30
       (.I0(data[5]),
        .O(modv_reg_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_31
       (.I0(data[0]),
        .O(modv_reg_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_32
       (.I0(data[4]),
        .O(modv_reg_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_33
       (.I0(data[3]),
        .O(modv_reg_i_33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_34
       (.I0(data[2]),
        .O(modv_reg_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    modv_reg_i_35
       (.I0(data[1]),
        .O(modv_reg_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_4
       (.I0(psin0[12]),
        .I1(phase),
        .I2(data[12]),
        .O(modv_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_5
       (.I0(psin0[11]),
        .I1(phase),
        .I2(data[11]),
        .O(modv_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_6
       (.I0(psin0[10]),
        .I1(phase),
        .I2(data[10]),
        .O(modv_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_7
       (.I0(psin0[9]),
        .I1(phase),
        .I2(data[9]),
        .O(modv_reg_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_8
       (.I0(psin0[8]),
        .I1(phase),
        .I2(data[8]),
        .O(modv_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    modv_reg_i_9
       (.I0(psin0[7]),
        .I1(phase),
        .I2(data[7]),
        .O(modv_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-12 {cell *THIS*}}" *) 
  DSP48E1 #(
    .ACASCREG(0),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(0),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(1),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    modvs_reg
       (.A({A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A[11],A}),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(\<const0>__0__0 ),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(reset),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({modvs_reg_n_58,modvs_reg_n_59,modvs_reg_n_60,modvs_reg_n_61,modvs_reg_n_62,modvs_reg_n_63,modvs_reg_n_64,modvs_reg_n_65,modvs_reg_n_66,modvs_reg_n_67,modvs_reg_n_68,modvs_reg_n_69,modvs_reg_n_70,modvs_reg_n_71,modvs_reg_n_72,modvs_reg_n_73,modvs_reg_n_74,modvs_reg_n_75,modvs_reg_n_76,modvs_reg_n_77,modvs_reg_n_78,modvs_reg_n_79,R,modvs_reg_n_96,modvs_reg_n_97,modvs_reg_n_98,modvs_reg_n_99,modvs_reg_n_100,modvs_reg_n_101,modvs_reg_n_102,modvs_reg_n_103,modvs_reg_n_104,modvs_reg_n_105}),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  DSP48E1 #(
    .ACASCREG(1),
    .ADREG(1),
    .ALUMODEREG(0),
    .AREG(1),
    .AUTORESET_PATDET("NO_RESET"),
    .A_INPUT("DIRECT"),
    .BCASCREG(0),
    .BREG(0),
    .B_INPUT("DIRECT"),
    .CARRYINREG(0),
    .CARRYINSELREG(0),
    .CREG(1),
    .DREG(1),
    .INMODEREG(0),
    .IS_ALUMODE_INVERTED(4'b0000),
    .IS_CARRYIN_INVERTED(1'b0),
    .IS_CLK_INVERTED(1'b0),
    .IS_INMODE_INVERTED(5'b00000),
    .IS_OPMODE_INVERTED(7'b0000000),
    .MASK(48'h3FFFFFFFFFFF),
    .MREG(1),
    .OPMODEREG(0),
    .PATTERN(48'h000000000000),
    .PREG(0),
    .SEL_MASK("MASK"),
    .SEL_PATTERN("PATTERN"),
    .USE_DPORT("FALSE"),
    .USE_MULT("MULTIPLY"),
    .USE_PATTERN_DETECT("NO_PATDET"),
    .USE_SIMD("ONE48")) 
    modys_reg
       (.A({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\I_6/output_reg_n_0_[10] ,\I_6/output_reg_n_0_[9] ,\I_6/output_reg_n_0_[8] ,\I_6/output_reg_n_0_[7] ,\I_6/output_reg_n_0_[6] ,\I_6/output_reg_n_0_[5] ,\I_6/output_reg_n_0_[4] ,\I_6/output_reg_n_0_[3] ,\I_6/output_reg_n_0_[2] ,\I_6/output_reg_n_0_[1] ,\I_6/output_reg_n_0_ }),
        .ACIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .ALUMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .B({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .BCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .C({VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2,VCC_2}),
        .CARRYCASCIN(\<const0>__0__0 ),
        .CARRYIN(\<const0>__0__0 ),
        .CARRYINSEL({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CEA1(\<const0>__0__0 ),
        .CEA2(reset),
        .CEAD(\<const0>__0__0 ),
        .CEALUMODE(\<const0>__0__0 ),
        .CEB1(\<const0>__0__0 ),
        .CEB2(\<const0>__0__0 ),
        .CEC(\<const0>__0__0 ),
        .CECARRYIN(\<const0>__0__0 ),
        .CECTRL(\<const0>__0__0 ),
        .CED(\<const0>__0__0 ),
        .CEINMODE(\<const0>__0__0 ),
        .CEM(reset),
        .CEP(\<const0>__0__0 ),
        .CLK(clk),
        .D({GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2,GND_2}),
        .INMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .MULTSIGNIN(\<const0>__0__0 ),
        .OPMODE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .P({modys_reg_n_58,modys_reg_n_59,modys_reg_n_60,modys_reg_n_61,modys_reg_n_62,modys_reg_n_63,modys_reg_n_64,modys_reg_n_65,modys_reg_n_66,modys_reg_n_67,modys_reg_n_68,modys_reg_n_69,modys_reg_n_70,modys_reg_n_71,modys_reg_n_72,modys_reg_n_73,modys_reg_n_74,modys_reg_n_75,modys_reg_n_76,modys_reg_n_77,modys_reg_n_78,modys_reg_n_79,modys_reg_n_80,modys_reg_n_81,modys_reg_n_82,modys_reg_n_83,modys_reg_n_84,modys_reg_n_85,modys_reg_n_86,modys_reg_n_87,modys_reg_n_88,modys_reg_n_89,modys_reg_n_90,modys_reg_n_91,modys_reg_n_92,modys_reg_n_93,modys_reg_n_94,modys_reg_n_95,modys_reg_n_96,modys_reg_n_97,modys_reg_n_98,modys_reg_n_99,modys_reg_n_100,modys_reg_n_101,modys_reg_n_102,modys_reg_n_103,modys_reg_n_104,modys_reg_n_105}),
        .PCIN({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .RSTA(\<const0>__0__0 ),
        .RSTALLCARRYIN(\<const0>__0__0 ),
        .RSTALUMODE(\<const0>__0__0 ),
        .RSTB(\<const0>__0__0 ),
        .RSTC(\<const0>__0__0 ),
        .RSTCTRL(\<const0>__0__0 ),
        .RSTD(\<const0>__0__0 ),
        .RSTINMODE(\<const0>__0__0 ),
        .RSTM(\<const0>__0__0 ),
        .RSTP(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_1
       (.I0(\I_5/multOp_carry__1_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp__39_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_1__0
       (.I0(\I_4/multOp_carry__1_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp__39_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_2
       (.I0(\I_5/multOp_carry__1_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp__39_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_2__0
       (.I0(\I_4/multOp_carry__1_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp__39_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_3
       (.I0(\I_5/multOp_carry__0_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp__39_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_3__0
       (.I0(\I_4/multOp_carry__0_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp__39_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_4
       (.I0(\I_5/multOp_carry__0_n_5 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_4 ),
        .O(multOp__39_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__0_i_4__0
       (.I0(\I_4/multOp_carry__0_n_5 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_4 ),
        .O(multOp__39_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_5
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_5 ),
        .I1(\I_5/multOp_carry__1_n_6 ),
        .I2(\I_5/multOp_carry__1_n_5 ),
        .I3(\I_5/plusOp_inferred__6_carry__0_n_4 ),
        .O(multOp__39_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_5__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_5 ),
        .I1(\I_4/multOp_carry__1_n_6 ),
        .I2(\I_4/multOp_carry__1_n_5 ),
        .I3(\I_4/plusOp_inferred__6_carry__0_n_4 ),
        .O(multOp__39_carry__0_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_6
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_6 ),
        .I1(\I_5/multOp_carry__1_n_7 ),
        .I2(\I_5/multOp_carry__1_n_6 ),
        .I3(\I_5/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp__39_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_6__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_6 ),
        .I1(\I_4/multOp_carry__1_n_7 ),
        .I2(\I_4/multOp_carry__1_n_6 ),
        .I3(\I_4/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp__39_carry__0_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_7
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_7 ),
        .I1(\I_5/multOp_carry__0_n_4 ),
        .I2(\I_5/multOp_carry__1_n_7 ),
        .I3(\I_5/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp__39_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_7__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_7 ),
        .I1(\I_4/multOp_carry__0_n_4 ),
        .I2(\I_4/multOp_carry__1_n_7 ),
        .I3(\I_4/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp__39_carry__0_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_8
       (.I0(\I_5/plusOp_inferred__6_carry_n_4 ),
        .I1(\I_5/multOp_carry__0_n_5 ),
        .I2(\I_5/multOp_carry__0_n_4 ),
        .I3(\I_5/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp__39_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__0_i_8__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_4 ),
        .I1(\I_4/multOp_carry__0_n_5 ),
        .I2(\I_4/multOp_carry__0_n_4 ),
        .I3(\I_4/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp__39_carry__0_i_8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__1_i_1
       (.I0(\I_5/multOp_carry__2_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__1_i_1__0
       (.I0(\I_4/multOp_carry__2_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__1_i_2
       (.I0(\I_5/multOp_carry__2_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp__39_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry__1_i_2__0
       (.I0(\I_4/multOp_carry__2_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp__39_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    multOp__39_carry__1_i_3
       (.I0(\I_5/multOp_carry__1_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .O(multOp__39_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    multOp__39_carry__1_i_3__0
       (.I0(\I_4/multOp_carry__1_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .O(multOp__39_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp__39_carry__1_i_4
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_5/multOp_carry__1_n_4 ),
        .O(multOp__39_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp__39_carry__1_i_4__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_4/multOp_carry__1_n_4 ),
        .O(multOp__39_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4BB4)) 
    multOp__39_carry__1_i_5
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_5 ),
        .I1(\I_5/multOp_carry__2_n_6 ),
        .I2(\I_5/multOp_carry__2_n_1 ),
        .I3(\I_5/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp__39_carry__1_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4BB4)) 
    multOp__39_carry__1_i_5__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_5 ),
        .I1(\I_4/multOp_carry__2_n_6 ),
        .I2(\I_4/multOp_carry__2_n_1 ),
        .I3(\I_4/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp__39_carry__1_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__1_i_6
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_6 ),
        .I1(\I_5/multOp_carry__2_n_7 ),
        .I2(\I_5/multOp_carry__2_n_6 ),
        .I3(\I_5/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry__1_i_6__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_6 ),
        .I1(\I_4/multOp_carry__2_n_7 ),
        .I2(\I_4/multOp_carry__2_n_6 ),
        .I3(\I_4/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    multOp__39_carry__1_i_7
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_5/multOp_carry__1_n_4 ),
        .I2(\I_5/multOp_carry__2_n_7 ),
        .I3(\I_5/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp__39_carry__1_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    multOp__39_carry__1_i_7__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_4/multOp_carry__1_n_4 ),
        .I2(\I_4/multOp_carry__2_n_7 ),
        .I3(\I_4/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp__39_carry__1_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6966)) 
    multOp__39_carry__1_i_8
       (.I0(\I_5/multOp_carry__1_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .I2(\I_5/plusOp_inferred__6_carry__0_n_4 ),
        .I3(\I_5/multOp_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6966)) 
    multOp__39_carry__1_i_8__0
       (.I0(\I_4/multOp_carry__1_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .I2(\I_4/plusOp_inferred__6_carry__0_n_4 ),
        .I3(\I_4/multOp_carry__1_n_5 ),
        .O(multOp__39_carry__1_i_8__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    multOp__39_carry__2_i_1
       (.I0(\I_5/multOp_carry__2_n_1 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp__39_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    multOp__39_carry__2_i_1__0
       (.I0(\I_4/multOp_carry__2_n_1 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp__39_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry_i_1
       (.I0(\I_5/multOp_carry__0_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_5 ),
        .O(multOp__39_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry_i_1__0
       (.I0(\I_4/multOp_carry__0_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_5 ),
        .O(multOp__39_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry_i_2
       (.I0(\I_5/multOp_carry__0_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_6 ),
        .O(multOp__39_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    multOp__39_carry_i_2__0
       (.I0(\I_4/multOp_carry__0_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_6 ),
        .O(multOp__39_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    multOp__39_carry_i_3
       (.I0(\I_5/multOp_carry_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_7 ),
        .O(multOp__39_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    multOp__39_carry_i_3__0
       (.I0(\I_4/multOp_carry_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_7 ),
        .O(multOp__39_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry_i_4
       (.I0(\I_5/plusOp_inferred__6_carry_n_5 ),
        .I1(\I_5/multOp_carry__0_n_6 ),
        .I2(\I_5/multOp_carry__0_n_5 ),
        .I3(\I_5/plusOp_inferred__6_carry_n_4 ),
        .O(multOp__39_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry_i_4__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_5 ),
        .I1(\I_4/multOp_carry__0_n_6 ),
        .I2(\I_4/multOp_carry__0_n_5 ),
        .I3(\I_4/plusOp_inferred__6_carry_n_4 ),
        .O(multOp__39_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry_i_5
       (.I0(\I_5/plusOp_inferred__6_carry_n_6 ),
        .I1(\I_5/multOp_carry__0_n_7 ),
        .I2(\I_5/multOp_carry__0_n_6 ),
        .I3(\I_5/plusOp_inferred__6_carry_n_5 ),
        .O(multOp__39_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB44B)) 
    multOp__39_carry_i_5__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_6 ),
        .I1(\I_4/multOp_carry__0_n_7 ),
        .I2(\I_4/multOp_carry__0_n_6 ),
        .I3(\I_4/plusOp_inferred__6_carry_n_5 ),
        .O(multOp__39_carry_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    multOp__39_carry_i_6
       (.I0(\I_5/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_5/multOp_carry_n_4 ),
        .I2(\I_5/multOp_carry__0_n_7 ),
        .I3(\I_5/plusOp_inferred__6_carry_n_6 ),
        .O(multOp__39_carry_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2DD2)) 
    multOp__39_carry_i_6__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_4/multOp_carry_n_4 ),
        .I2(\I_4/multOp_carry__0_n_7 ),
        .I3(\I_4/plusOp_inferred__6_carry_n_6 ),
        .O(multOp__39_carry_i_6__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp__39_carry_i_7
       (.I0(\I_5/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_5/multOp_carry_n_4 ),
        .O(multOp__39_carry_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp__39_carry_i_7__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_4/multOp_carry_n_4 ),
        .O(multOp__39_carry_i_7__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_1
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_4 ),
        .O(multOp_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_1__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_4 ),
        .O(multOp_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_2
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_2__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_5 ),
        .O(multOp_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_3
       (.I0(\I_5/plusOp_inferred__6_carry_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_3__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_6 ),
        .O(multOp_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_4
       (.I0(\I_5/plusOp_inferred__6_carry_n_5 ),
        .I1(\I_5/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__0_i_4__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_5 ),
        .I1(\I_4/plusOp_inferred__6_carry__0_n_7 ),
        .O(multOp_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp_carry__1_i_1
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    multOp_carry__1_i_1__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_2
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_2__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_3
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_4 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_3__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_4 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_6 ),
        .O(multOp_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_4
       (.I0(\I_5/plusOp_inferred__6_carry__0_n_5 ),
        .I1(\I_5/plusOp_inferred__6_carry__1_n_7 ),
        .O(multOp_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry__1_i_4__0
       (.I0(\I_4/plusOp_inferred__6_carry__0_n_5 ),
        .I1(\I_4/plusOp_inferred__6_carry__1_n_7 ),
        .O(multOp_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry__2_i_1
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry__2_i_1__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_4 ),
        .O(multOp_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry__2_i_2
       (.I0(\I_5/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry__2_i_2__0
       (.I0(\I_4/plusOp_inferred__6_carry__1_n_5 ),
        .O(multOp_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry_i_1
       (.I0(\I_5/plusOp_inferred__6_carry_n_6 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_4 ),
        .O(multOp_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry_i_1__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_6 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_4 ),
        .O(multOp_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry_i_2
       (.I0(\I_5/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_5/plusOp_inferred__6_carry_n_5 ),
        .O(multOp_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    multOp_carry_i_2__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_7 ),
        .I1(\I_4/plusOp_inferred__6_carry_n_5 ),
        .O(multOp_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry_i_3
       (.I0(\I_5/plusOp_inferred__6_carry_n_6 ),
        .O(multOp_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    multOp_carry_i_3__0
       (.I0(\I_4/plusOp_inferred__6_carry_n_6 ),
        .O(multOp_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h002A80AA)) 
    \output[0]_i_1 
       (.I0(sync),
        .I1(en_bild),
        .I2(tmr_austastung),
        .I3(\output_reg[0]_i_2_n_7 ),
        .I4(plusOp0_in[0]),
        .O(\output[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_10 
       (.I0(\output_reg[0]_i_2_n_6 ),
        .I1(modys_reg_n_94),
        .O(\output[0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_11 
       (.I0(\output_reg[0]_i_2_n_7 ),
        .I1(modys_reg_n_95),
        .O(\output[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_4 
       (.I0(L[3]),
        .I1(R[3]),
        .O(\output[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_5 
       (.I0(L[2]),
        .I1(R[2]),
        .O(\output[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_6 
       (.I0(L[1]),
        .I1(R[1]),
        .O(\output[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_7 
       (.I0(L[0]),
        .I1(R[0]),
        .O(\output[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_8 
       (.I0(\output_reg[0]_i_2_n_4 ),
        .I1(modys_reg_n_92),
        .O(\output[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[0]_i_9 
       (.I0(\output_reg[0]_i_2_n_5 ),
        .I1(modys_reg_n_93),
        .O(\output[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[10]_i_1 
       (.I0(sync),
        .I1(\output_reg[12]_i_2_n_6 ),
        .O(\output[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[11]_i_1 
       (.I0(sync),
        .I1(\output_reg[12]_i_2_n_5 ),
        .O(\output[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[12]_i_1 
       (.I0(sync),
        .I1(\output_reg[12]_i_2_n_4 ),
        .O(\output[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_10 
       (.I0(\output_reg[12]_i_8_n_5 ),
        .I1(modys_reg_n_85),
        .O(\output[12]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_11 
       (.I0(\output_reg[12]_i_8_n_6 ),
        .I1(modys_reg_n_86),
        .O(\output[12]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_12 
       (.I0(\output_reg[12]_i_8_n_7 ),
        .I1(modys_reg_n_87),
        .O(\output[12]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_13 
       (.I0(L[11]),
        .I1(R[11]),
        .O(\output[12]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_14 
       (.I0(L[10]),
        .I1(R[10]),
        .O(\output[12]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_15 
       (.I0(L[9]),
        .I1(R[9]),
        .O(\output[12]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_16 
       (.I0(L[8]),
        .I1(R[8]),
        .O(\output[12]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[12]_i_3 
       (.I0(plusOp0_in[12]),
        .I1(\output_reg[15]_i_8_n_7 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[12]_i_4 
       (.I0(plusOp0_in[11]),
        .I1(\output_reg[12]_i_8_n_4 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[12]_i_5 
       (.I0(plusOp0_in[10]),
        .I1(\output_reg[12]_i_8_n_5 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[12]_i_6 
       (.I0(plusOp0_in[9]),
        .I1(\output_reg[12]_i_8_n_6 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[12]_i_9 
       (.I0(\output_reg[12]_i_8_n_4 ),
        .I1(modys_reg_n_84),
        .O(\output[12]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[13]_i_1 
       (.I0(sync),
        .I1(\output_reg[15]_i_3_n_7 ),
        .O(\output[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[14]_i_1 
       (.I0(sync),
        .I1(\output_reg[15]_i_3_n_6 ),
        .O(\output[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[15]_i_1 
       (.I0(sync),
        .I1(\output_reg[15]_i_3_n_5 ),
        .O(\output[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_10 
       (.I0(\output_reg[15]_i_8_n_5 ),
        .I1(modys_reg_n_81),
        .O(\output[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_11 
       (.I0(\output_reg[15]_i_8_n_6 ),
        .I1(modys_reg_n_82),
        .O(\output[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_12 
       (.I0(\output_reg[15]_i_8_n_7 ),
        .I1(modys_reg_n_83),
        .O(\output[15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_13 
       (.I0(L[15]),
        .I1(R[15]),
        .O(\output[15]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_14 
       (.I0(L[14]),
        .I1(R[14]),
        .O(\output[15]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_15 
       (.I0(L[13]),
        .I1(R[13]),
        .O(\output[15]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_16 
       (.I0(L[12]),
        .I1(R[12]),
        .O(\output[15]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \output[15]_i_2 
       (.I0(reset),
        .O(clear));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[15]_i_4 
       (.I0(plusOp0_in[15]),
        .I1(\output_reg[15]_i_8_n_4 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[15]_i_5 
       (.I0(plusOp0_in[14]),
        .I1(\output_reg[15]_i_8_n_5 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[15]_i_6 
       (.I0(plusOp0_in[13]),
        .I1(\output_reg[15]_i_8_n_6 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[15]_i_9 
       (.I0(\output_reg[15]_i_8_n_4 ),
        .I1(modys_reg_n_80),
        .O(\output[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[1]_i_1 
       (.I0(sync),
        .I1(\output_reg[4]_i_2_n_7 ),
        .O(\output[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[2]_i_1 
       (.I0(sync),
        .I1(\output_reg[4]_i_2_n_6 ),
        .O(\output[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[3]_i_1 
       (.I0(sync),
        .I1(\output_reg[4]_i_2_n_5 ),
        .O(\output[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[4]_i_1 
       (.I0(sync),
        .I1(\output_reg[4]_i_2_n_4 ),
        .O(\output[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[4]_i_3 
       (.I0(plusOp0_in[0]),
        .I1(\output_reg[0]_i_2_n_7 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[4]_i_4 
       (.I0(plusOp0_in[4]),
        .I1(\output_reg[8]_i_8_n_7 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[4]_i_5 
       (.I0(plusOp0_in[3]),
        .I1(\output_reg[0]_i_2_n_4 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[4]_i_6 
       (.I0(plusOp0_in[2]),
        .I1(\output_reg[0]_i_2_n_5 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[4]_i_7 
       (.I0(plusOp0_in[1]),
        .I1(\output_reg[0]_i_2_n_6 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[5]_i_1 
       (.I0(sync),
        .I1(\output_reg[8]_i_2_n_7 ),
        .O(\output[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[6]_i_1 
       (.I0(sync),
        .I1(\output_reg[8]_i_2_n_6 ),
        .O(\output[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[7]_i_1 
       (.I0(sync),
        .I1(\output_reg[8]_i_2_n_5 ),
        .O(\output[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[8]_i_1 
       (.I0(sync),
        .I1(\output_reg[8]_i_2_n_4 ),
        .O(\output[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_10 
       (.I0(\output_reg[8]_i_8_n_5 ),
        .I1(modys_reg_n_89),
        .O(\output[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_11 
       (.I0(\output_reg[8]_i_8_n_6 ),
        .I1(modys_reg_n_90),
        .O(\output[8]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_12 
       (.I0(\output_reg[8]_i_8_n_7 ),
        .I1(modys_reg_n_91),
        .O(\output[8]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_13 
       (.I0(L[7]),
        .I1(R[7]),
        .O(\output[8]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_14 
       (.I0(L[6]),
        .I1(R[6]),
        .O(\output[8]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_15 
       (.I0(L[5]),
        .I1(R[5]),
        .O(\output[8]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_16 
       (.I0(L[4]),
        .I1(R[4]),
        .O(\output[8]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hACCC)) 
    \output[8]_i_3 
       (.I0(plusOp0_in[8]),
        .I1(\output_reg[12]_i_8_n_7 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(prevideo[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[8]_i_4 
       (.I0(plusOp0_in[7]),
        .I1(\output_reg[8]_i_8_n_4 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[8]_i_5 
       (.I0(plusOp0_in[6]),
        .I1(\output_reg[8]_i_8_n_5 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5333)) 
    \output[8]_i_6 
       (.I0(plusOp0_in[5]),
        .I1(\output_reg[8]_i_8_n_6 ),
        .I2(tmr_austastung),
        .I3(en_bild),
        .O(\output[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \output[8]_i_9 
       (.I0(\output_reg[8]_i_8_n_4 ),
        .I1(modys_reg_n_88),
        .O(\output[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \output[9]_i_1 
       (.I0(sync),
        .I1(\output_reg[12]_i_2_n_7 ),
        .O(\output[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[0]_i_1_n_0 ),
        .Q(\output [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[0]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO(output_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[3:0]),
        .O({\output_reg[0]_i_2_n_4 ,\output_reg[0]_i_2_n_5 ,\output_reg[0]_i_2_n_6 ,\output_reg[0]_i_2_n_7 }),
        .S({\output[0]_i_4_n_0 ,\output[0]_i_5_n_0 ,\output[0]_i_6_n_0 ,\output[0]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[0]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\output_reg[0]_i_3_n_0 ,\output_reg[0]_i_3_n_1 ,\output_reg[0]_i_3_n_2 ,\output_reg[0]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\output_reg[0]_i_2_n_4 ,\output_reg[0]_i_2_n_5 ,\output_reg[0]_i_2_n_6 ,\output_reg[0]_i_2_n_7 }),
        .O(plusOp0_in[3:0]),
        .S({\output[0]_i_8_n_0 ,\output[0]_i_9_n_0 ,\output[0]_i_10_n_0 ,\output[0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[10]_i_1_n_0 ),
        .Q(\output [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[11]_i_1_n_0 ),
        .Q(\output [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[12]_i_1_n_0 ),
        .Q(\output [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[12]_i_2 
       (.CI(\output_reg[8]_i_2_n_0 ),
        .CO({\output_reg[12]_i_2_n_0 ,\output_reg[12]_i_2_n_1 ,\output_reg[12]_i_2_n_2 ,\output_reg[12]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\output_reg[12]_i_2_n_4 ,\output_reg[12]_i_2_n_5 ,\output_reg[12]_i_2_n_6 ,\output_reg[12]_i_2_n_7 }),
        .S({\output[12]_i_3_n_0 ,\output[12]_i_4_n_0 ,prevideo[10:9]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[12]_i_7 
       (.CI(\output_reg[8]_i_7_n_0 ),
        .CO({\output_reg[12]_i_7_n_0 ,\output_reg[12]_i_7_n_1 ,\output_reg[12]_i_7_n_2 ,\output_reg[12]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\output_reg[12]_i_8_n_4 ,\output_reg[12]_i_8_n_5 ,\output_reg[12]_i_8_n_6 ,\output_reg[12]_i_8_n_7 }),
        .O(plusOp0_in[11:8]),
        .S({\output[12]_i_9_n_0 ,\output[12]_i_10_n_0 ,\output[12]_i_11_n_0 ,\output[12]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[12]_i_8 
       (.CI(\output_reg[8]_i_8_n_0 ),
        .CO({\output_reg[12]_i_8_n_0 ,\output_reg[12]_i_8_n_1 ,\output_reg[12]_i_8_n_2 ,\output_reg[12]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[11:8]),
        .O({\output_reg[12]_i_8_n_4 ,\output_reg[12]_i_8_n_5 ,\output_reg[12]_i_8_n_6 ,\output_reg[12]_i_8_n_7 }),
        .S({\output[12]_i_13_n_0 ,\output[12]_i_14_n_0 ,\output[12]_i_15_n_0 ,\output[12]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[13]_i_1_n_0 ),
        .Q(\output [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[14]_i_1_n_0 ),
        .Q(\output [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[15]_i_1_n_0 ),
        .Q(\output [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[15]_i_3 
       (.CI(\output_reg[12]_i_2_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\output_reg[15]_i_3_n_4 ,\output_reg[15]_i_3_n_5 ,\output_reg[15]_i_3_n_6 ,\output_reg[15]_i_3_n_7 }),
        .S({\<const0>__0__0 ,prevideo[15:14],\output[15]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[15]_i_7 
       (.CI(\output_reg[12]_i_7_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\output_reg[15]_i_8_n_5 ,\output_reg[15]_i_8_n_6 ,\output_reg[15]_i_8_n_7 }),
        .O(plusOp0_in[15:12]),
        .S({\output[15]_i_9_n_0 ,\output[15]_i_10_n_0 ,\output[15]_i_11_n_0 ,\output[15]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[15]_i_8 
       (.CI(\output_reg[12]_i_8_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,L[14:12]}),
        .O({\output_reg[15]_i_8_n_4 ,\output_reg[15]_i_8_n_5 ,\output_reg[15]_i_8_n_6 ,\output_reg[15]_i_8_n_7 }),
        .S({\output[15]_i_13_n_0 ,\output[15]_i_14_n_0 ,\output[15]_i_15_n_0 ,\output[15]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[1]_i_1_n_0 ),
        .Q(\output [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[2]_i_1_n_0 ),
        .Q(\output [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[3]_i_1_n_0 ),
        .Q(\output [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[4]_i_1_n_0 ),
        .Q(\output [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[4]_i_2 
       (.CI(\<const0>__0__0 ),
        .CO({\output_reg[4]_i_2_n_0 ,\output_reg[4]_i_2_n_1 ,\output_reg[4]_i_2_n_2 ,\output_reg[4]_i_2_n_3 }),
        .CYINIT(prevideo[0]),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 }),
        .O({\output_reg[4]_i_2_n_4 ,\output_reg[4]_i_2_n_5 ,\output_reg[4]_i_2_n_6 ,\output_reg[4]_i_2_n_7 }),
        .S({prevideo[4:2],\output[4]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[5]_i_1_n_0 ),
        .Q(\output [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[6]_i_1_n_0 ),
        .Q(\output [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[7]_i_1_n_0 ),
        .Q(\output [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[8]_i_1_n_0 ),
        .Q(\output [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[8]_i_2 
       (.CI(\output_reg[4]_i_2_n_0 ),
        .CO({\output_reg[8]_i_2_n_0 ,\output_reg[8]_i_2_n_1 ,\output_reg[8]_i_2_n_2 ,\output_reg[8]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\output_reg[8]_i_2_n_4 ,\output_reg[8]_i_2_n_5 ,\output_reg[8]_i_2_n_6 ,\output_reg[8]_i_2_n_7 }),
        .S({prevideo[8],\output[8]_i_4_n_0 ,\output[8]_i_5_n_0 ,\output[8]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[8]_i_7 
       (.CI(\output_reg[0]_i_3_n_0 ),
        .CO({\output_reg[8]_i_7_n_0 ,\output_reg[8]_i_7_n_1 ,\output_reg[8]_i_7_n_2 ,\output_reg[8]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\output_reg[8]_i_8_n_4 ,\output_reg[8]_i_8_n_5 ,\output_reg[8]_i_8_n_6 ,\output_reg[8]_i_8_n_7 }),
        .O(plusOp0_in[7:4]),
        .S({\output[8]_i_9_n_0 ,\output[8]_i_10_n_0 ,\output[8]_i_11_n_0 ,\output[8]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \output_reg[8]_i_8 
       (.CI(output_reg[3]),
        .CO({\output_reg[8]_i_8_n_0 ,\output_reg[8]_i_8_n_1 ,\output_reg[8]_i_8_n_2 ,\output_reg[8]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(L[7:4]),
        .O({\output_reg[8]_i_8_n_4 ,\output_reg[8]_i_8_n_5 ,\output_reg[8]_i_8_n_6 ,\output_reg[8]_i_8_n_7 }),
        .S({\output[8]_i_13_n_0 ,\output[8]_i_14_n_0 ,\output[8]_i_15_n_0 ,\output[8]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \output_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .CLR(clear),
        .D(\output[9]_i_1_n_0 ),
        .Q(\output [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__0_i_1
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr2_carry__4_n_5 ),
        .I2(\I_0/pixctr2_carry__4_n_7 ),
        .O(pixctr1_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__0_i_2
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr2_carry__3_n_4 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(pixctr1_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__0_i_3
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr2_carry__3_n_7 ),
        .I2(\I_0/pixctr2_carry__2_n_5 ),
        .O(pixctr1_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__0_i_4
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr2_carry__2_n_6 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(pixctr1_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    pixctr1_carry__1_i_1
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .O(pixctr1_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__1_i_2
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr2_carry__6_n_7 ),
        .I2(\I_0/pixctr2_carry__5_n_5 ),
        .O(pixctr1_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry__1_i_3
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr2_carry__5_n_6 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(pixctr1_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    pixctr1_carry_i_1
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr2_carry__1_n_7 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(pixctr1_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    pixctr1_carry_i_2
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr2_carry__0_n_5 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(pixctr1_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    pixctr1_carry_i_3
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .I2(\I_0/pixctr2_carry_n_5 ),
        .O(pixctr1_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    pixctr1_carry_i_4
       (.I0(\I_0/pixctr2_carry_n_6 ),
        .I1(\I_0/pixctr_reg_n_0_ ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(pixctr1_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \pixctr[0]_i_1 
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[10]_i_1 
       (.I0(\I_0/pixctr2_carry__1_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[11]_i_1 
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[12]_i_1 
       (.I0(\I_0/pixctr2_carry__1_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[13]_i_1 
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[14]_i_1 
       (.I0(\I_0/pixctr2_carry__2_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[15]_i_1 
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[16]_i_1 
       (.I0(\I_0/pixctr2_carry__2_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[17]_i_1 
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[18]_i_1 
       (.I0(\I_0/pixctr2_carry__3_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[19]_i_1 
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[1]_i_1 
       (.I0(\I_0/pixctr2_carry_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[20]_i_1 
       (.I0(\I_0/pixctr2_carry__3_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[21]_i_1 
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[22]_i_1 
       (.I0(\I_0/pixctr2_carry__4_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[23]_i_1 
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[24]_i_1 
       (.I0(\I_0/pixctr2_carry__4_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[25]_i_1 
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[26]_i_1 
       (.I0(\I_0/pixctr2_carry__5_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[27]_i_1 
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[28]_i_1 
       (.I0(\I_0/pixctr2_carry__5_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[29]_i_1 
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[2]_i_1 
       (.I0(\I_0/pixctr2_carry_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[30]_i_1 
       (.I0(\I_0/pixctr2_carry__6_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[31]_i_1 
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \pixctr[31]_i_2 
       (.I0(reset),
        .O(pixctr));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[3]_i_1 
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[4]_i_1 
       (.I0(\I_0/pixctr2_carry_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[5]_i_1 
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[6]_i_1 
       (.I0(\I_0/pixctr2_carry__0_n_6 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[7]_i_1 
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[8]_i_1 
       (.I0(\I_0/pixctr2_carry__0_n_4 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \pixctr[9]_i_1 
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(\I_0/pixctr [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry__0_i_1
       (.I0(g0_b6_n_0),
        .I1(g0_b6__0_n_0),
        .I2(g0_b6__1_n_0),
        .O(plusOp__0_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair4" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry__0_i_2
       (.I0(g0_b5_n_0),
        .I1(g0_b5__0_n_0),
        .I2(g0_b5__1_n_0),
        .O(plusOp__0_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair3" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry__0_i_3
       (.I0(g0_b4_n_0),
        .I1(g0_b4__0_n_0),
        .I2(g0_b4__1_n_0),
        .O(plusOp__0_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair2" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry__0_i_4
       (.I0(g0_b3_n_0),
        .I1(g0_b3__0_n_0),
        .I2(g0_b3__1_n_0),
        .O(plusOp__0_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hE81717E8)) 
    plusOp__0_carry__0_i_5
       (.I0(g0_b6__1_n_0),
        .I1(g0_b6__0_n_0),
        .I2(g0_b6_n_0),
        .I3(g0_b7_n_0),
        .I4(g0_b7__0_n_0),
        .O(plusOp__0_carry__0_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry__0_i_6
       (.I0(plusOp__0_carry__0_i_2_n_0),
        .I1(g0_b6__0_n_0),
        .I2(g0_b6_n_0),
        .I3(g0_b6__1_n_0),
        .O(plusOp__0_carry__0_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair4" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry__0_i_7
       (.I0(g0_b5_n_0),
        .I1(g0_b5__0_n_0),
        .I2(g0_b5__1_n_0),
        .I3(plusOp__0_carry__0_i_3_n_0),
        .O(plusOp__0_carry__0_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair3" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry__0_i_8
       (.I0(g0_b4_n_0),
        .I1(g0_b4__0_n_0),
        .I2(g0_b4__1_n_0),
        .I3(plusOp__0_carry__0_i_4_n_0),
        .O(plusOp__0_carry__0_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    plusOp__0_carry__1_i_1
       (.I0(g0_b7_n_0),
        .I1(g0_b7__0_n_0),
        .O(plusOp__0_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8778)) 
    plusOp__0_carry__1_i_2
       (.I0(g0_b7__0_n_0),
        .I1(g0_b7_n_0),
        .I2(g0_b8_n_0),
        .I3(g0_b8__0_n_0),
        .O(plusOp__0_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair1" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry_i_1
       (.I0(g0_b2_n_0),
        .I1(g0_b2__0_n_0),
        .I2(g0_b2__1_n_0),
        .O(plusOp__0_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair0" *) 
  LUT3 #(
    .INIT(8'hE8)) 
    plusOp__0_carry_i_2
       (.I0(g0_b1_n_0),
        .I1(g0_b1__0_n_0),
        .I2(g0_b1__1_n_0),
        .O(plusOp__0_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair2" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry_i_3
       (.I0(g0_b3_n_0),
        .I1(g0_b3__0_n_0),
        .I2(g0_b3__1_n_0),
        .I3(plusOp__0_carry_i_1_n_0),
        .O(plusOp__0_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair1" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry_i_4
       (.I0(g0_b2_n_0),
        .I1(g0_b2__0_n_0),
        .I2(g0_b2__1_n_0),
        .I3(plusOp__0_carry_i_2_n_0),
        .O(plusOp__0_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* HLUTNM = "lutpair0" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    plusOp__0_carry_i_5
       (.I0(g0_b1_n_0),
        .I1(g0_b1__0_n_0),
        .I2(g0_b1__1_n_0),
        .I3(g0_b0__0_n_0),
        .O(plusOp__0_carry_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8F800000707FFFFF))
    plusOp_inferred__3_carry__0_i_1
       (.I0(\I_3/multOp_n_88 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\I_5/sr_reg_n_0_[14][7] ),
        .O(plusOp_inferred__3_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__0_i_1__0
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp__0_n_88 ),
        .I3(en_bild),
        .I4(\sr_reg[14] [7]),
        .O(plusOp_inferred__3_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__0_i_2
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_89 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][6] ),
        .O(plusOp_inferred__3_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__0_i_2__0
       (.I0(\I_3/multOp__0_n_89 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [6]),
        .O(plusOp_inferred__3_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__0_i_3
       (.I0(\I_3/multOp_n_90 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\I_5/sr_reg_n_0_[14][5] ),
        .O(plusOp_inferred__3_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__0_i_3__0
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp__0_n_90 ),
        .I3(en_bild),
        .I4(\sr_reg[14] [5]),
        .O(plusOp_inferred__3_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__0_i_4
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_91 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][4] ),
        .O(plusOp_inferred__3_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__0_i_4__0
       (.I0(\I_3/multOp__0_n_91 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [4]),
        .O(plusOp_inferred__3_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__1_i_1
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_84 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][11] ),
        .O(plusOp_inferred__3_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__1_i_1__0
       (.I0(\I_3/multOp__0_n_84 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [11]),
        .O(plusOp_inferred__3_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__1_i_2
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_85 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][10] ),
        .O(plusOp_inferred__3_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__1_i_2__0
       (.I0(\I_3/multOp__0_n_85 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [10]),
        .O(plusOp_inferred__3_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__1_i_3
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_86 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][9] ),
        .O(plusOp_inferred__3_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__1_i_3__0
       (.I0(\I_3/multOp__0_n_86 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [9]),
        .O(plusOp_inferred__3_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry__1_i_4
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_87 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][8] ),
        .O(plusOp_inferred__3_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry__1_i_4__0
       (.I0(\I_3/multOp__0_n_87 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [8]),
        .O(plusOp_inferred__3_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry_i_1
       (.I0(\I_3/multOp_n_92 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\I_5/sr_reg_n_0_[14][3] ),
        .O(plusOp_inferred__3_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry_i_1__0
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp__0_n_92 ),
        .I3(en_bild),
        .I4(\sr_reg[14] [3]),
        .O(plusOp_inferred__3_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry_i_2
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp_n_93 ),
        .I3(en_bild),
        .I4(\I_5/sr_reg_n_0_[14][2] ),
        .O(plusOp_inferred__3_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry_i_2__0
       (.I0(\I_3/multOp__0_n_93 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [2]),
        .O(plusOp_inferred__3_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry_i_3
       (.I0(\I_3/multOp_n_94 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\I_5/sr_reg_n_0_[14][1] ),
        .O(plusOp_inferred__3_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFF8000)) 
    plusOp_inferred__3_carry_i_3__0
       (.I0(tmr_austastung),
        .I1(sr_reg),
        .I2(\I_3/multOp__0_n_94 ),
        .I3(en_bild),
        .I4(\sr_reg[14] [1]),
        .O(plusOp_inferred__3_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry_i_4
       (.I0(\I_3/multOp_n_95 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\I_5/sr_reg_n_0_[14][0] ),
        .O(plusOp_inferred__3_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h707FFFFF8F800000)) 
    plusOp_inferred__3_carry_i_4__0
       (.I0(\I_3/multOp__0_n_95 ),
        .I1(sr_reg),
        .I2(en_bild),
        .I3(tmr_en_burst),
        .I4(tmr_austastung),
        .I5(\sr_reg[14] [0]),
        .O(plusOp_inferred__3_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_1
       (.I0(\I_5/sr_reg_n_0_[1][7] ),
        .I1(\I_5/sr_reg_n_0_[12][7] ),
        .O(plusOp_inferred__5_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_1__0
       (.I0(\sr_reg[1] [7]),
        .I1(\sr_reg[12] [7]),
        .O(plusOp_inferred__5_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_2
       (.I0(\I_5/sr_reg_n_0_[1][6] ),
        .I1(\I_5/sr_reg_n_0_[12][6] ),
        .O(plusOp_inferred__5_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_2__0
       (.I0(\sr_reg[1] [6]),
        .I1(\sr_reg[12] [6]),
        .O(plusOp_inferred__5_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_3
       (.I0(\I_5/sr_reg_n_0_[1][5] ),
        .I1(\I_5/sr_reg_n_0_[12][5] ),
        .O(plusOp_inferred__5_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_3__0
       (.I0(\sr_reg[1] [5]),
        .I1(\sr_reg[12] [5]),
        .O(plusOp_inferred__5_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_4
       (.I0(\I_5/sr_reg_n_0_[1][4] ),
        .I1(\I_5/sr_reg_n_0_[12][4] ),
        .O(plusOp_inferred__5_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__0_i_4__0
       (.I0(\sr_reg[1] [4]),
        .I1(\sr_reg[12] [4]),
        .O(plusOp_inferred__5_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_1
       (.I0(\I_5/sr_reg_n_0_[1][11] ),
        .I1(\I_5/sr_reg_n_0_[12][11] ),
        .O(plusOp_inferred__5_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_1__0
       (.I0(\sr_reg[1] [11]),
        .I1(\sr_reg[12] [11]),
        .O(plusOp_inferred__5_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_2
       (.I0(\I_5/sr_reg_n_0_[1][10] ),
        .I1(\I_5/sr_reg_n_0_[12][10] ),
        .O(plusOp_inferred__5_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_2__0
       (.I0(\sr_reg[1] [10]),
        .I1(\sr_reg[12] [10]),
        .O(plusOp_inferred__5_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_3
       (.I0(\I_5/sr_reg_n_0_[1][9] ),
        .I1(\I_5/sr_reg_n_0_[12][9] ),
        .O(plusOp_inferred__5_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_3__0
       (.I0(\sr_reg[1] [9]),
        .I1(\sr_reg[12] [9]),
        .O(plusOp_inferred__5_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_4
       (.I0(\I_5/sr_reg_n_0_[1][8] ),
        .I1(\I_5/sr_reg_n_0_[12][8] ),
        .O(plusOp_inferred__5_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry__1_i_4__0
       (.I0(\sr_reg[1] [8]),
        .I1(\sr_reg[12] [8]),
        .O(plusOp_inferred__5_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_1
       (.I0(\I_5/sr_reg_n_0_[1][3] ),
        .I1(\I_5/sr_reg_n_0_[12][3] ),
        .O(plusOp_inferred__5_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_1__0
       (.I0(\sr_reg[1] [3]),
        .I1(\sr_reg[12] [3]),
        .O(plusOp_inferred__5_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_2
       (.I0(\I_5/sr_reg_n_0_[1][2] ),
        .I1(\I_5/sr_reg_n_0_[12][2] ),
        .O(plusOp_inferred__5_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_2__0
       (.I0(\sr_reg[1] [2]),
        .I1(\sr_reg[12] [2]),
        .O(plusOp_inferred__5_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_3
       (.I0(\I_5/sr_reg_n_0_[1][1] ),
        .I1(\I_5/sr_reg_n_0_[12][1] ),
        .O(plusOp_inferred__5_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_3__0
       (.I0(\sr_reg[1] [1]),
        .I1(\sr_reg[12] [1]),
        .O(plusOp_inferred__5_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_4
       (.I0(\I_5/sr_reg_n_0_[1][0] ),
        .I1(\I_5/sr_reg_n_0_[12][0] ),
        .O(plusOp_inferred__5_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__5_carry_i_4__0
       (.I0(\sr_reg[1] [0]),
        .I1(\sr_reg[12] [0]),
        .O(plusOp_inferred__5_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_1
       (.I0(\I_5/sr_reg_n_0_[0][7] ),
        .I1(\I_5/sr_reg_n_0_[13][7] ),
        .O(plusOp_inferred__6_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_1__0
       (.I0(\sr_reg[0] [7]),
        .I1(\sr_reg[13] [7]),
        .O(plusOp_inferred__6_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_2
       (.I0(\I_5/sr_reg_n_0_[0][6] ),
        .I1(\I_5/sr_reg_n_0_[13][6] ),
        .O(plusOp_inferred__6_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_2__0
       (.I0(\sr_reg[0] [6]),
        .I1(\sr_reg[13] [6]),
        .O(plusOp_inferred__6_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_3
       (.I0(\I_5/sr_reg_n_0_[0][5] ),
        .I1(\I_5/sr_reg_n_0_[13][5] ),
        .O(plusOp_inferred__6_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_3__0
       (.I0(\sr_reg[0] [5]),
        .I1(\sr_reg[13] [5]),
        .O(plusOp_inferred__6_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_4
       (.I0(\I_5/sr_reg_n_0_[0][4] ),
        .I1(\I_5/sr_reg_n_0_[13][4] ),
        .O(plusOp_inferred__6_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__0_i_4__0
       (.I0(\sr_reg[0] [4]),
        .I1(\sr_reg[13] [4]),
        .O(plusOp_inferred__6_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_1
       (.I0(\I_5/sr_reg_n_0_[0][11] ),
        .I1(\I_5/sr_reg_n_0_[13][11] ),
        .O(plusOp_inferred__6_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_1__0
       (.I0(\sr_reg[0] [11]),
        .I1(\sr_reg[13] [11]),
        .O(plusOp_inferred__6_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_2
       (.I0(\I_5/sr_reg_n_0_[0][10] ),
        .I1(\I_5/sr_reg_n_0_[13][10] ),
        .O(plusOp_inferred__6_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_2__0
       (.I0(\sr_reg[0] [10]),
        .I1(\sr_reg[13] [10]),
        .O(plusOp_inferred__6_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_3
       (.I0(\I_5/sr_reg_n_0_[0][9] ),
        .I1(\I_5/sr_reg_n_0_[13][9] ),
        .O(plusOp_inferred__6_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_3__0
       (.I0(\sr_reg[0] [9]),
        .I1(\sr_reg[13] [9]),
        .O(plusOp_inferred__6_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_4
       (.I0(\I_5/sr_reg_n_0_[0][8] ),
        .I1(\I_5/sr_reg_n_0_[13][8] ),
        .O(plusOp_inferred__6_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry__1_i_4__0
       (.I0(\sr_reg[0] [8]),
        .I1(\sr_reg[13] [8]),
        .O(plusOp_inferred__6_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_1
       (.I0(\I_5/sr_reg_n_0_[0][3] ),
        .I1(\I_5/sr_reg_n_0_[13][3] ),
        .O(plusOp_inferred__6_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_1__0
       (.I0(\sr_reg[0] [3]),
        .I1(\sr_reg[13] [3]),
        .O(plusOp_inferred__6_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_2
       (.I0(\I_5/sr_reg_n_0_[0][2] ),
        .I1(\I_5/sr_reg_n_0_[13][2] ),
        .O(plusOp_inferred__6_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_2__0
       (.I0(\sr_reg[0] [2]),
        .I1(\sr_reg[13] [2]),
        .O(plusOp_inferred__6_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_3
       (.I0(\I_5/sr_reg_n_0_[0][1] ),
        .I1(\I_5/sr_reg_n_0_[13][1] ),
        .O(plusOp_inferred__6_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_3__0
       (.I0(\sr_reg[0] [1]),
        .I1(\sr_reg[13] [1]),
        .O(plusOp_inferred__6_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_4
       (.I0(\I_5/sr_reg_n_0_ ),
        .I1(\I_5/sr_reg_n_0_[13][0] ),
        .O(plusOp_inferred__6_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__6_carry_i_4__0
       (.I0(\sr_reg[0] [0]),
        .I1(\sr_reg[13] [0]),
        .O(plusOp_inferred__6_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_1
       (.I0(\I_5/multOp__39_carry__0_n_7 ),
        .I1(C[7]),
        .O(plusOp_inferred__7__62_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_1__0
       (.I0(multOp0[7]),
        .I1(C__0[7]),
        .O(plusOp_inferred__7__62_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_2
       (.I0(\I_5/multOp__39_carry_n_4 ),
        .I1(C[6]),
        .O(plusOp_inferred__7__62_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_2__0
       (.I0(multOp0[6]),
        .I1(C__0[6]),
        .O(plusOp_inferred__7__62_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_3
       (.I0(\I_5/multOp__39_carry_n_5 ),
        .I1(C[5]),
        .O(plusOp_inferred__7__62_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_3__0
       (.I0(multOp0[5]),
        .I1(C__0[5]),
        .O(plusOp_inferred__7__62_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_4
       (.I0(\I_5/multOp__39_carry_n_6 ),
        .I1(C[4]),
        .O(plusOp_inferred__7__62_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__0_i_4__0
       (.I0(multOp0[4]),
        .I1(C__0[4]),
        .O(plusOp_inferred__7__62_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_1
       (.I0(\I_5/multOp__39_carry__1_n_7 ),
        .I1(C[11]),
        .O(plusOp_inferred__7__62_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_1__0
       (.I0(multOp0[11]),
        .I1(C__0[11]),
        .O(plusOp_inferred__7__62_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_2
       (.I0(\I_5/multOp__39_carry__0_n_4 ),
        .I1(C[10]),
        .O(plusOp_inferred__7__62_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_2__0
       (.I0(multOp0[10]),
        .I1(C__0[10]),
        .O(plusOp_inferred__7__62_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_3
       (.I0(\I_5/multOp__39_carry__0_n_5 ),
        .I1(C[9]),
        .O(plusOp_inferred__7__62_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_3__0
       (.I0(multOp0[9]),
        .I1(C__0[9]),
        .O(plusOp_inferred__7__62_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_4
       (.I0(\I_5/multOp__39_carry__0_n_6 ),
        .I1(C[8]),
        .O(plusOp_inferred__7__62_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__1_i_4__0
       (.I0(multOp0[8]),
        .I1(C__0[8]),
        .O(plusOp_inferred__7__62_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    plusOp_inferred__7__62_carry__2_i_1
       (.I0(C[15]),
        .O(plusOp_inferred__7__62_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    plusOp_inferred__7__62_carry__2_i_1__0
       (.I0(C__0[15]),
        .O(plusOp_inferred__7__62_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_2
       (.I0(C[15]),
        .I1(\I_5/multOp__39_carry__2_n_7 ),
        .O(plusOp_inferred__7__62_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_2__0
       (.I0(C__0[15]),
        .I1(multOp0[15]),
        .O(plusOp_inferred__7__62_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_3
       (.I0(\I_5/multOp__39_carry__1_n_4 ),
        .I1(C[14]),
        .O(plusOp_inferred__7__62_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_3__0
       (.I0(multOp0[14]),
        .I1(C__0[14]),
        .O(plusOp_inferred__7__62_carry__2_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_4
       (.I0(\I_5/multOp__39_carry__1_n_5 ),
        .I1(C[13]),
        .O(plusOp_inferred__7__62_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_4__0
       (.I0(multOp0[13]),
        .I1(C__0[13]),
        .O(plusOp_inferred__7__62_carry__2_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_5
       (.I0(\I_5/multOp__39_carry__1_n_6 ),
        .I1(C[12]),
        .O(plusOp_inferred__7__62_carry__2_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry__2_i_5__0
       (.I0(multOp0[12]),
        .I1(C__0[12]),
        .O(plusOp_inferred__7__62_carry__2_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_1
       (.I0(C[18]),
        .I1(C[19]),
        .O(plusOp_inferred__7__62_carry__3_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_1__0
       (.I0(C__0[18]),
        .I1(C__0[19]),
        .O(plusOp_inferred__7__62_carry__3_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_2
       (.I0(C[17]),
        .I1(C[18]),
        .O(plusOp_inferred__7__62_carry__3_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_2__0
       (.I0(C__0[17]),
        .I1(C__0[18]),
        .O(plusOp_inferred__7__62_carry__3_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_3
       (.I0(C[16]),
        .I1(C[17]),
        .O(plusOp_inferred__7__62_carry__3_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_3__0
       (.I0(C__0[16]),
        .I1(C__0[17]),
        .O(plusOp_inferred__7__62_carry__3_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_4
       (.I0(C[15]),
        .I1(C[16]),
        .O(plusOp_inferred__7__62_carry__3_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__3_i_4__0
       (.I0(C__0[15]),
        .I1(C__0[16]),
        .O(plusOp_inferred__7__62_carry__3_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_1
       (.I0(C[21]),
        .I1(C[22]),
        .O(plusOp_inferred__7__62_carry__4_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_1__0
       (.I0(C__0[21]),
        .I1(C__0[22]),
        .O(plusOp_inferred__7__62_carry__4_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_2
       (.I0(C[20]),
        .I1(C[21]),
        .O(plusOp_inferred__7__62_carry__4_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_2__0
       (.I0(C__0[20]),
        .I1(C__0[21]),
        .O(plusOp_inferred__7__62_carry__4_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_3
       (.I0(C[19]),
        .I1(C[20]),
        .O(plusOp_inferred__7__62_carry__4_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7__62_carry__4_i_3__0
       (.I0(C__0[19]),
        .I1(C__0[20]),
        .O(plusOp_inferred__7__62_carry__4_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_1
       (.I0(\I_5/multOp__39_carry_n_7 ),
        .I1(C[3]),
        .O(plusOp_inferred__7__62_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_1__0
       (.I0(multOp0[3]),
        .I1(C__0[3]),
        .O(plusOp_inferred__7__62_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_2
       (.I0(\I_5/multOp_carry_n_5 ),
        .I1(C[2]),
        .O(plusOp_inferred__7__62_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_2__0
       (.I0(multOp0[2]),
        .I1(C__0[2]),
        .O(plusOp_inferred__7__62_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_3
       (.I0(\I_5/multOp_carry_n_6 ),
        .I1(C[1]),
        .O(plusOp_inferred__7__62_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_3__0
       (.I0(multOp0[1]),
        .I1(C__0[1]),
        .O(plusOp_inferred__7__62_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_4
       (.I0(\I_5/multOp_carry_n_7 ),
        .I1(\I_5/plusOp__3_n_105 ),
        .O(plusOp_inferred__7__62_carry_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7__62_carry_i_4__0
       (.I0(multOp0[0]),
        .I1(\I_4/plusOp__3_n_105 ),
        .O(plusOp_inferred__7__62_carry_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_1
       (.I0(\I_5/multOp__0 [6]),
        .I1(\I_5/plusOp__3_n_97 ),
        .O(plusOp_inferred__7_carry__0_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_1__0
       (.I0(\I_4/multOp__0 [6]),
        .I1(\I_4/plusOp__3_n_97 ),
        .O(plusOp_inferred__7_carry__0_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_2
       (.I0(\I_5/multOp__0 [5]),
        .I1(\I_5/plusOp__3_n_98 ),
        .O(plusOp_inferred__7_carry__0_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_2__0
       (.I0(\I_4/multOp__0 [5]),
        .I1(\I_4/plusOp__3_n_98 ),
        .O(plusOp_inferred__7_carry__0_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_3
       (.I0(\I_5/multOp__0 [4]),
        .I1(\I_5/plusOp__3_n_99 ),
        .O(plusOp_inferred__7_carry__0_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_3__0
       (.I0(\I_4/multOp__0 [4]),
        .I1(\I_4/plusOp__3_n_99 ),
        .O(plusOp_inferred__7_carry__0_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_4
       (.I0(\I_5/multOp__0 [3]),
        .I1(\I_5/plusOp__3_n_100 ),
        .O(plusOp_inferred__7_carry__0_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__0_i_4__0
       (.I0(\I_4/multOp__0 [3]),
        .I1(\I_4/plusOp__3_n_100 ),
        .O(plusOp_inferred__7_carry__0_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_1
       (.I0(\I_5/multOp__0 [10]),
        .I1(\I_5/plusOp__3_n_93 ),
        .O(plusOp_inferred__7_carry__1_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_1__0
       (.I0(\I_4/multOp__0 [10]),
        .I1(\I_4/plusOp__3_n_93 ),
        .O(plusOp_inferred__7_carry__1_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_2
       (.I0(\I_5/multOp__0 [9]),
        .I1(\I_5/plusOp__3_n_94 ),
        .O(plusOp_inferred__7_carry__1_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_2__0
       (.I0(\I_4/multOp__0 [9]),
        .I1(\I_4/plusOp__3_n_94 ),
        .O(plusOp_inferred__7_carry__1_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_3
       (.I0(\I_5/multOp__0 [8]),
        .I1(\I_5/plusOp__3_n_95 ),
        .O(plusOp_inferred__7_carry__1_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_3__0
       (.I0(\I_4/multOp__0 [8]),
        .I1(\I_4/plusOp__3_n_95 ),
        .O(plusOp_inferred__7_carry__1_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_4
       (.I0(\I_5/multOp__0 [7]),
        .I1(\I_5/plusOp__3_n_96 ),
        .O(plusOp_inferred__7_carry__1_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__1_i_4__0
       (.I0(\I_4/multOp__0 [7]),
        .I1(\I_4/plusOp__3_n_96 ),
        .O(plusOp_inferred__7_carry__1_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    plusOp_inferred__7_carry__2_i_1
       (.I0(\I_5/plusOp__3_n_92 ),
        .O(plusOp_inferred__7_carry__2_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    plusOp_inferred__7_carry__2_i_1__0
       (.I0(\I_4/plusOp__3_n_92 ),
        .O(plusOp_inferred__7_carry__2_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_2
       (.I0(\I_5/plusOp__3_n_90 ),
        .I1(\I_5/plusOp__3_n_89 ),
        .O(plusOp_inferred__7_carry__2_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_2__0
       (.I0(\I_4/plusOp__3_n_90 ),
        .I1(\I_4/plusOp__3_n_89 ),
        .O(plusOp_inferred__7_carry__2_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_3
       (.I0(\I_5/plusOp__3_n_91 ),
        .I1(\I_5/plusOp__3_n_90 ),
        .O(plusOp_inferred__7_carry__2_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_3__0
       (.I0(\I_4/plusOp__3_n_91 ),
        .I1(\I_4/plusOp__3_n_90 ),
        .O(plusOp_inferred__7_carry__2_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_4
       (.I0(\I_5/plusOp__3_n_92 ),
        .I1(\I_5/plusOp__3_n_91 ),
        .O(plusOp_inferred__7_carry__2_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__2_i_4__0
       (.I0(\I_4/plusOp__3_n_92 ),
        .I1(\I_4/plusOp__3_n_91 ),
        .O(plusOp_inferred__7_carry__2_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__2_i_5
       (.I0(\I_5/plusOp__3_n_92 ),
        .I1(\I_5/multOp__0 [11]),
        .O(plusOp_inferred__7_carry__2_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry__2_i_5__0
       (.I0(\I_4/plusOp__3_n_92 ),
        .I1(\I_4/multOp__0 [11]),
        .O(plusOp_inferred__7_carry__2_i_5__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_1
       (.I0(\I_5/plusOp__3_n_86 ),
        .I1(\I_5/plusOp__3_n_85 ),
        .O(plusOp_inferred__7_carry__3_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_1__0
       (.I0(\I_4/plusOp__3_n_86 ),
        .I1(\I_4/plusOp__3_n_85 ),
        .O(plusOp_inferred__7_carry__3_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_2
       (.I0(\I_5/plusOp__3_n_87 ),
        .I1(\I_5/plusOp__3_n_86 ),
        .O(plusOp_inferred__7_carry__3_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_2__0
       (.I0(\I_4/plusOp__3_n_87 ),
        .I1(\I_4/plusOp__3_n_86 ),
        .O(plusOp_inferred__7_carry__3_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_3
       (.I0(\I_5/plusOp__3_n_88 ),
        .I1(\I_5/plusOp__3_n_87 ),
        .O(plusOp_inferred__7_carry__3_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_3__0
       (.I0(\I_4/plusOp__3_n_88 ),
        .I1(\I_4/plusOp__3_n_87 ),
        .O(plusOp_inferred__7_carry__3_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_4
       (.I0(\I_5/plusOp__3_n_89 ),
        .I1(\I_5/plusOp__3_n_88 ),
        .O(plusOp_inferred__7_carry__3_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__3_i_4__0
       (.I0(\I_4/plusOp__3_n_89 ),
        .I1(\I_4/plusOp__3_n_88 ),
        .O(plusOp_inferred__7_carry__3_i_4__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__4_i_1
       (.I0(\I_5/plusOp__3_n_84 ),
        .I1(\I_5/plusOp__3_n_83 ),
        .O(plusOp_inferred__7_carry__4_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__4_i_1__0
       (.I0(\I_4/plusOp__3_n_84 ),
        .I1(\I_4/plusOp__3_n_83 ),
        .O(plusOp_inferred__7_carry__4_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__4_i_2
       (.I0(\I_5/plusOp__3_n_85 ),
        .I1(\I_5/plusOp__3_n_84 ),
        .O(plusOp_inferred__7_carry__4_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    plusOp_inferred__7_carry__4_i_2__0
       (.I0(\I_4/plusOp__3_n_85 ),
        .I1(\I_4/plusOp__3_n_84 ),
        .O(plusOp_inferred__7_carry__4_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_1
       (.I0(\I_5/multOp__0 [2]),
        .I1(\I_5/plusOp__3_n_101 ),
        .O(plusOp_inferred__7_carry_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_1__0
       (.I0(\I_4/multOp__0 [2]),
        .I1(\I_4/plusOp__3_n_101 ),
        .O(plusOp_inferred__7_carry_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_2
       (.I0(\I_5/multOp__0 [1]),
        .I1(\I_5/plusOp__3_n_102 ),
        .O(plusOp_inferred__7_carry_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_2__0
       (.I0(\I_4/multOp__0 [1]),
        .I1(\I_4/plusOp__3_n_102 ),
        .O(plusOp_inferred__7_carry_i_2__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_3
       (.I0(\I_5/multOp__0 [0]),
        .I1(\I_5/plusOp__3_n_103 ),
        .O(plusOp_inferred__7_carry_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    plusOp_inferred__7_carry_i_3__0
       (.I0(\I_4/multOp__0 [0]),
        .I1(\I_4/plusOp__3_n_103 ),
        .O(plusOp_inferred__7_carry_i_3__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][0]_i_1 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp_n_95 ),
        .O(pre_yuv_v[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][0]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_95 ),
        .O(\input [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][10]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_85 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][10]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_85 ),
        .O(\input [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][11]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_84 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][11]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_84 ),
        .O(\input [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][1]_i_1 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp_n_94 ),
        .O(pre_yuv_v[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][1]_i_1__0 
       (.I0(en_bild),
        .I1(\I_3/multOp__0_n_94 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(\input [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][2]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_93 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][2]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_93 ),
        .O(\input [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][3]_i_1 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp_n_92 ),
        .O(pre_yuv_v[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][3]_i_1__0 
       (.I0(en_bild),
        .I1(\I_3/multOp__0_n_92 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(\input [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][4]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_91 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][4]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_91 ),
        .O(\input [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][5]_i_1 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp_n_90 ),
        .O(pre_yuv_v[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][5]_i_1__0 
       (.I0(en_bild),
        .I1(\I_3/multOp__0_n_90 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(\input [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][6]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_89 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][6]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_89 ),
        .O(\input [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][7]_i_1 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp_n_88 ),
        .O(pre_yuv_v[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][7]_i_1__0 
       (.I0(en_bild),
        .I1(\I_3/multOp__0_n_88 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(\input [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sr[0][7]_i_2 
       (.I0(reset),
        .O(sr));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][8]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_87 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][8]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_87 ),
        .O(\input [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \sr[0][9]_i_1 
       (.I0(en_bild),
        .I1(\I_3/multOp_n_86 ),
        .I2(sr_reg),
        .I3(tmr_austastung),
        .O(pre_yuv_v[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA8080808)) 
    \sr[0][9]_i_1__0 
       (.I0(tmr_austastung),
        .I1(tmr_en_burst),
        .I2(en_bild),
        .I3(sr_reg),
        .I4(\I_3/multOp__0_n_86 ),
        .O(\input [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \sr[2][7]_i_1 
       (.I0(reset),
        .O(\sr[2][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDCE #(
    .INIT(1'b0),
    .IS_CLR_INVERTED(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0)) 
    \sr_reg[0][11]_i_2 
       (.C(clk15M),
        .CE(\<const1>__0__0 ),
        .CLR(sr),
        .D(\<const1>__0__0 ),
        .Q(sr_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1DDDFFFF1DDD3333)) 
    sync_i_1
       (.I0(sync_i_2_n_0),
        .I1(i_sync_c),
        .I2(\I_0/i_phase433_in ),
        .I3(\I_0/i_phase4 ),
        .I4(\i_sync_c[1]_i_1_n_0 ),
        .I5(sync_i_3_n_0),
        .O(\I_0/p_1_in ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_10
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(sync_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_11
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(sync_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    sync_i_13
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(sync_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    sync_i_14
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(sync_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_15
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(sync_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_16
       (.I0(\I_0/pixctr2_carry__5_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_6 ),
        .O(sync_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_17
       (.I0(\I_0/pixctr2_carry__5_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_4 ),
        .O(sync_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_19
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(sync_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF888)) 
    sync_i_2
       (.I0(\I_0/i_en_verteq2 ),
        .I1(\I_0/i_phase4 ),
        .I2(\I_0/i_en_verteq1 ),
        .I3(\I_0/i_en_vertbr1 ),
        .O(sync_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_20
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(sync_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_21
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(sync_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_22
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(sync_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_24
       (.I0(\I_0/pixctr2_carry__4_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__4_n_6 ),
        .O(sync_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_25
       (.I0(\I_0/pixctr2_carry__4_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_4 ),
        .O(sync_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_26
       (.I0(\I_0/pixctr2_carry__3_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__3_n_6 ),
        .O(sync_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_27
       (.I0(\I_0/pixctr2_carry__3_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_4 ),
        .O(sync_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_29
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(sync_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0777)) 
    sync_i_3
       (.I0(\I_0/i_en_vertbr1 ),
        .I1(\I_0/i_en_vertbr131_in ),
        .I2(\I_0/i_en_vertbr2 ),
        .I3(\I_0/i_phase4 ),
        .O(sync_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_30
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(sync_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_31
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(sync_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_32
       (.I0(\I_0/pixctr2_carry__1_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(sync_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    sync_i_34
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__1_n_7 ),
        .O(sync_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_35
       (.I0(\I_0/pixctr2_carry__2_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__2_n_6 ),
        .O(sync_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_36
       (.I0(\I_0/pixctr2_carry__2_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_4 ),
        .O(sync_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_37
       (.I0(\I_0/pixctr2_carry__1_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__1_n_6 ),
        .O(sync_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    sync_i_38
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__1_n_7 ),
        .I2(\I_0/pixctr2_carry__0_n_4 ),
        .O(sync_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    sync_i_39
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .O(sync_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    sync_i_40
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_7 ),
        .O(sync_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_41
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(sync_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    sync_i_42
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__0_n_7 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(sync_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_43
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(sync_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    sync_i_44
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(sync_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    sync_i_45
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry_n_7 ),
        .O(sync_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_46
       (.I0(\I_0/pixctr2_carry__0_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__0_n_6 ),
        .O(sync_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_47
       (.I0(\I_0/pixctr2_carry__0_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_4 ),
        .O(sync_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_48
       (.I0(\I_0/pixctr2_carry_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_6 ),
        .O(sync_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    sync_i_49
       (.I0(\I_0/pixctr_reg_n_0_ ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry_n_7 ),
        .O(sync_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    sync_i_7
       (.I0(\I_0/pixctr2_carry__6_n_5 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .O(sync_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    sync_i_8
       (.I0(\I_0/pixctr1_carry__1_n_1 ),
        .I1(\I_0/pixctr2_carry__6_n_6 ),
        .I2(\I_0/pixctr2_carry__6_n_5 ),
        .O(sync_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCD)) 
    sync_i_9
       (.I0(\I_0/pixctr2_carry__6_n_7 ),
        .I1(\I_0/pixctr1_carry__1_n_1 ),
        .I2(\I_0/pixctr2_carry__5_n_4 ),
        .O(sync_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_12
       (.CI(sync_reg_i_23_n_0),
        .CO({sync_reg_i_12_n_0,sync_reg_i_12_n_1,sync_reg_i_12_n_2,sync_reg_i_12_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({sync_i_24_n_0,sync_i_25_n_0,sync_i_26_n_0,sync_i_27_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_18
       (.CI(sync_reg_i_28_n_0),
        .CO({sync_reg_i_18_n_0,sync_reg_i_18_n_1,sync_reg_i_18_n_2,sync_reg_i_18_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({sync_i_29_n_0,sync_i_30_n_0,sync_i_31_n_0,sync_i_32_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_23
       (.CI(sync_reg_i_33_n_0),
        .CO({sync_reg_i_23_n_0,sync_reg_i_23_n_1,sync_reg_i_23_n_2,sync_reg_i_23_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,sync_i_34_n_0}),
        .S({sync_i_35_n_0,sync_i_36_n_0,sync_i_37_n_0,sync_i_38_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_28
       (.CI(\<const0>__0__0 ),
        .CO({sync_reg_i_28_n_0,sync_reg_i_28_n_1,sync_reg_i_28_n_2,sync_reg_i_28_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,sync_i_39_n_0,\<const0>__0__0 ,sync_i_40_n_0}),
        .S({sync_i_41_n_0,sync_i_42_n_0,sync_i_43_n_0,sync_i_44_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_33
       (.CI(\<const0>__0__0 ),
        .CO({sync_reg_i_33_n_0,sync_reg_i_33_n_1,sync_reg_i_33_n_2,sync_reg_i_33_n_3}),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,sync_i_45_n_0}),
        .S({sync_i_46_n_0,sync_i_47_n_0,sync_i_48_n_0,sync_i_49_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_4
       (.CI(sync_reg_i_6_n_0),
        .CO({\I_0/i_en_verteq2 ,sync_reg_i_4_n_1,sync_reg_i_4_n_2,sync_reg_i_4_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({sync_i_7_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({sync_i_8_n_0,sync_i_9_n_0,sync_i_10_n_0,sync_i_11_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_5
       (.CI(sync_reg_i_12_n_0),
        .CO({\I_0/i_en_verteq1 ,sync_reg_i_5_n_1,sync_reg_i_5_n_2,sync_reg_i_5_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({sync_i_13_n_0,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({sync_i_14_n_0,sync_i_15_n_0,sync_i_16_n_0,sync_i_17_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 sync_reg_i_6
       (.CI(sync_reg_i_18_n_0),
        .CO({sync_reg_i_6_n_0,sync_reg_i_6_n_1,sync_reg_i_6_n_2,sync_reg_i_6_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({sync_i_19_n_0,sync_i_20_n_0,sync_i_21_n_0,sync_i_22_n_0}));
endmodule
