module counter(input clk_i, rst_i, en_i, output blink_o);
endmodule // counter