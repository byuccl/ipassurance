module irqmp
   (rst,
    clk,
    .\apbi[psel] ({apbi[0],apbi[1],apbi[2],apbi[3],apbi[4],apbi[5],apbi[6],apbi[7],apbi[8],apbi[9],apbi[10],apbi[11],apbi[12],apbi[13],apbi[14],apbi[15]}),
    \apbi[penable] ,
    \apbi[paddr] ,
    \apbi[pwrite] ,
    \apbi[pwdata] ,
    \apbi[pirq] ,
    \apbi[testen] ,
    \apbi[testrst] ,
    \apbi[scanen] ,
    \apbi[testoen] ,
    \apbi[testin] ,
    \apbo[prdata] ,
    \apbo[pirq] ,
    \apbo[pconfig][0] ,
    \apbo[pconfig][1] ,
    \apbo[pindex] ,
    .\irqi[0][intack] (irqi),
    \irqi[0][irl] ,
    \irqi[0][pwd] ,
    \irqi[0][fpen] ,
    \irqi[0][err] ,
    \irqi[1][intack] ,
    \irqi[1][irl] ,
    \irqi[1][pwd] ,
    \irqi[1][fpen] ,
    \irqi[1][err] ,
    \irqi[2][intack] ,
    \irqi[2][irl] ,
    \irqi[2][pwd] ,
    \irqi[2][fpen] ,
    \irqi[2][err] ,
    \irqi[3][intack] ,
    \irqi[3][irl] ,
    \irqi[3][pwd] ,
    \irqi[3][fpen] ,
    \irqi[3][err] ,
    \irqo[0][irl] ,
    \irqo[0][resume] ,
    \irqo[0][rstrun] ,
    \irqo[0][rstvec] ,
    \irqo[0][index] ,
    \irqo[0][pwdsetaddr] ,
    \irqo[0][pwdnewaddr] ,
    \irqo[0][forceerr] ,
    \irqo[0][svtclrtt] ,
    \irqo[1][irl] ,
    \irqo[1][resume] ,
    \irqo[1][rstrun] ,
    \irqo[1][rstvec] ,
    \irqo[1][index] ,
    \irqo[1][pwdsetaddr] ,
    \irqo[1][pwdnewaddr] ,
    \irqo[1][forceerr] ,
    \irqo[1][svtclrtt] ,
    \irqo[2][irl] ,
    \irqo[2][resume] ,
    \irqo[2][rstrun] ,
    \irqo[2][rstvec] ,
    \irqo[2][index] ,
    \irqo[2][pwdsetaddr] ,
    \irqo[2][pwdnewaddr] ,
    \irqo[2][forceerr] ,
    \irqo[2][svtclrtt] ,
    \irqo[3][irl] ,
    \irqo[3][resume] ,
    \irqo[3][rstrun] ,
    \irqo[3][rstvec] ,
    \irqo[3][index] ,
    \irqo[3][pwdsetaddr] ,
    \irqo[3][pwdnewaddr] ,
    \irqo[3][forceerr] ,
    \irqo[3][svtclrtt] );
  input rst;
  input clk;
  input \apbi[penable] ;
  input [31:0]\apbi[paddr] ;
  input \apbi[pwrite] ;
  input [31:0]\apbi[pwdata] ;
  input [31:0]\apbi[pirq] ;
  input \apbi[testen] ;
  input \apbi[testrst] ;
  input \apbi[scanen] ;
  input \apbi[testoen] ;
  input [3:0]\apbi[testin] ;
  output [31:0]\apbo[prdata] ;
  output [31:0]\apbo[pirq] ;
  output [31:0]\apbo[pconfig][0] ;
  output [31:0]\apbo[pconfig][1] ;
  output [3:0]\apbo[pindex] ;
  input [3:0]\irqi[0][irl] ;
  input \irqi[0][pwd] ;
  input \irqi[0][fpen] ;
  input \irqi[0][err] ;
  input \irqi[1][intack] ;
  input [3:0]\irqi[1][irl] ;
  input \irqi[1][pwd] ;
  input \irqi[1][fpen] ;
  input \irqi[1][err] ;
  input \irqi[2][intack] ;
  input [3:0]\irqi[2][irl] ;
  input \irqi[2][pwd] ;
  input \irqi[2][fpen] ;
  input \irqi[2][err] ;
  input \irqi[3][intack] ;
  input [3:0]\irqi[3][irl] ;
  input \irqi[3][pwd] ;
  input \irqi[3][fpen] ;
  input \irqi[3][err] ;
  output [3:0]\irqo[0][irl] ;
  output \irqo[0][resume] ;
  output \irqo[0][rstrun] ;
  output [31:12]\irqo[0][rstvec] ;
  output [3:0]\irqo[0][index] ;
  output \irqo[0][pwdsetaddr] ;
  output [31:2]\irqo[0][pwdnewaddr] ;
  output \irqo[0][forceerr] ;
  output \irqo[0][svtclrtt] ;
  output [3:0]\irqo[1][irl] ;
  output \irqo[1][resume] ;
  output \irqo[1][rstrun] ;
  output [31:12]\irqo[1][rstvec] ;
  output [3:0]\irqo[1][index] ;
  output \irqo[1][pwdsetaddr] ;
  output [31:2]\irqo[1][pwdnewaddr] ;
  output \irqo[1][forceerr] ;
  output \irqo[1][svtclrtt] ;
  output [3:0]\irqo[2][irl] ;
  output \irqo[2][resume] ;
  output \irqo[2][rstrun] ;
  output [31:12]\irqo[2][rstvec] ;
  output [3:0]\irqo[2][index] ;
  output \irqo[2][pwdsetaddr] ;
  output [31:2]\irqo[2][pwdnewaddr] ;
  output \irqo[2][forceerr] ;
  output \irqo[2][svtclrtt] ;
  output [3:0]\irqo[3][irl] ;
  output \irqo[3][resume] ;
  output \irqo[3][rstrun] ;
  output [31:12]\irqo[3][rstvec] ;
  output [3:0]\irqo[3][index] ;
  output \irqo[3][pwdsetaddr] ;
  output [31:2]\irqo[3][pwdnewaddr] ;
  output \irqo[3][forceerr] ;
  output \irqo[3][svtclrtt] ;
  input [0:15]apbi;
  input irqi;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:15]apbi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbi[paddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbi[penable] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbi[pirq] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\apbi[pwdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbi[pwrite] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire apbo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [26:0]\^apbo[prdata] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][0]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][10]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][11]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][12]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][13]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][14]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][15]_INST_0_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][1]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][2]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][3]_INST_0_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][4]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][5]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][6]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][7]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][8]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \apbo[prdata][9]_INST_0_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire irqi;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[0][err] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqi[0][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[0][pwd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[1][err] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[1][intack] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqi[1][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[1][pwd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[2][err] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[2][intack] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqi[2][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[2][pwd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[3][err] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[3][intack] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqi[3][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqi[3][pwd] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire irqo;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[0][forceerr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqo[0][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[0][resume] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[0][svtclrtt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[1][forceerr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqo[1][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[1][resume] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[1][svtclrtt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[2][forceerr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqo[2][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[2][resume] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[2][svtclrtt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[3][forceerr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:1]\^irqo[3][index] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\irqo[3][irl] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:2]\irqo[3][pwdnewaddr] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[3][resume] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \irqo[3][svtclrtt] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in10_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in12_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in14_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in16_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in18_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in20_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in22_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in24_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in26_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in28_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in30_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in4_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in6_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_in8_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:1]p_5_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [15:1]p_6_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[clkcount][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[clkcount][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[clkcount][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cpurst][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[cpurst][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[forceerr][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][0][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][1][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][2][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[iforce][3][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[imask][0][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[imask][1][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[imask][2][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[ipend][9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][0][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][1][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][2][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[irl][3][3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[newaddr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[newaddr][2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddr][0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddr][0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddr][1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddr][2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddr][3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r[setaddrboot]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[clkcount_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[clkcount_n_0_][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[ibroadcast_n_0_][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[iforce][0]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[iforce][1]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[iforce][2]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[iforce][3]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[imask][0]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[imask][1]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[imask][2]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [14:0]\r_reg[imask][3]__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_reg[setaddrboot_n_0_] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire v;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\v[cpurst]1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[ibroadcast] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[ilevel] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[imask][0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[imask][1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[imask][2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \v[imask][3] ;

  assign \apbo[pconfig][0] [31] = irqo;
  assign \apbo[pconfig][0] [30] = irqo;
  assign \apbo[pconfig][0] [29] = irqo;
  assign \apbo[pconfig][0] [28] = irqo;
  assign \apbo[pconfig][0] [27] = irqo;
  assign \apbo[pconfig][0] [26] = irqo;
  assign \apbo[pconfig][0] [25] = irqo;
  assign \apbo[pconfig][0] [24] = \^irqo[3][index] [1];
  assign \apbo[pconfig][0] [23] = irqo;
  assign \apbo[pconfig][0] [22] = irqo;
  assign \apbo[pconfig][0] [21] = irqo;
  assign \apbo[pconfig][0] [20] = irqo;
  assign \apbo[pconfig][0] [19] = irqo;
  assign \apbo[pconfig][0] [18] = irqo;
  assign \apbo[pconfig][0] [17] = irqo;
  assign \apbo[pconfig][0] [16] = irqo;
  assign \apbo[pconfig][0] [15] = \^irqo[3][index] [1];
  assign \apbo[pconfig][0] [14] = \^irqo[3][index] [1];
  assign \apbo[pconfig][0] [13] = irqo;
  assign \apbo[pconfig][0] [12] = \^irqo[3][index] [1];
  assign \apbo[pconfig][0] [11] = irqo;
  assign \apbo[pconfig][0] [10] = irqo;
  assign \apbo[pconfig][0] [9] = irqo;
  assign \apbo[pconfig][0] [8] = irqo;
  assign \apbo[pconfig][0] [7] = \^irqo[3][index] [1];
  assign \apbo[pconfig][0] [6] = irqo;
  assign \apbo[pconfig][0] [5] = irqo;
  assign \apbo[pconfig][0] [4] = irqo;
  assign \apbo[pconfig][0] [3] = irqo;
  assign \apbo[pconfig][0] [2] = irqo;
  assign \apbo[pconfig][0] [1] = irqo;
  assign \apbo[pconfig][0] [0] = irqo;
  assign \apbo[pconfig][1] [31] = irqo;
  assign \apbo[pconfig][1] [30] = irqo;
  assign \apbo[pconfig][1] [29] = irqo;
  assign \apbo[pconfig][1] [28] = irqo;
  assign \apbo[pconfig][1] [27] = irqo;
  assign \apbo[pconfig][1] [26] = irqo;
  assign \apbo[pconfig][1] [25] = irqo;
  assign \apbo[pconfig][1] [24] = irqo;
  assign \apbo[pconfig][1] [23] = irqo;
  assign \apbo[pconfig][1] [22] = irqo;
  assign \apbo[pconfig][1] [21] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [20] = irqo;
  assign \apbo[pconfig][1] [19] = irqo;
  assign \apbo[pconfig][1] [18] = irqo;
  assign \apbo[pconfig][1] [17] = irqo;
  assign \apbo[pconfig][1] [16] = irqo;
  assign \apbo[pconfig][1] [15] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [14] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [13] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [12] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [11] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [10] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [9] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [8] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [7] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [6] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [5] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [4] = \^irqo[3][index] [1];
  assign \apbo[pconfig][1] [3] = irqo;
  assign \apbo[pconfig][1] [2] = irqo;
  assign \apbo[pconfig][1] [1] = irqo;
  assign \apbo[pconfig][1] [0] = \^irqo[3][index] [1];
  assign \apbo[pindex] [3] = irqo;
  assign \apbo[pindex] [2] = irqo;
  assign \apbo[pindex] [1] = \^irqo[3][index] [1];
  assign \apbo[pindex] [0] = irqo;
  assign \apbo[pirq] [31] = irqo;
  assign \apbo[pirq] [30] = irqo;
  assign \apbo[pirq] [29] = irqo;
  assign \apbo[pirq] [28] = irqo;
  assign \apbo[pirq] [27] = irqo;
  assign \apbo[pirq] [26] = irqo;
  assign \apbo[pirq] [25] = irqo;
  assign \apbo[pirq] [24] = irqo;
  assign \apbo[pirq] [23] = irqo;
  assign \apbo[pirq] [22] = irqo;
  assign \apbo[pirq] [21] = irqo;
  assign \apbo[pirq] [20] = irqo;
  assign \apbo[pirq] [19] = irqo;
  assign \apbo[pirq] [18] = irqo;
  assign \apbo[pirq] [17] = irqo;
  assign \apbo[pirq] [16] = irqo;
  assign \apbo[pirq] [15] = irqo;
  assign \apbo[pirq] [14] = irqo;
  assign \apbo[pirq] [13] = irqo;
  assign \apbo[pirq] [12] = irqo;
  assign \apbo[pirq] [11] = irqo;
  assign \apbo[pirq] [10] = irqo;
  assign \apbo[pirq] [9] = irqo;
  assign \apbo[pirq] [8] = irqo;
  assign \apbo[pirq] [7] = irqo;
  assign \apbo[pirq] [6] = irqo;
  assign \apbo[pirq] [5] = irqo;
  assign \apbo[pirq] [4] = irqo;
  assign \apbo[pirq] [3] = irqo;
  assign \apbo[pirq] [2] = irqo;
  assign \apbo[pirq] [1] = irqo;
  assign \apbo[pirq] [0] = irqo;
  assign \apbo[prdata] [31] = irqo;
  assign \apbo[prdata] [30] = irqo;
  assign \apbo[prdata] [29] = apbo;
  assign \apbo[prdata] [28] = apbo;
  assign \apbo[prdata] [27] = apbo;
  assign \apbo[prdata] [26] = \^apbo[prdata] [26];
  assign \apbo[prdata] [25] = irqo;
  assign \apbo[prdata] [24] = irqo;
  assign \apbo[prdata] [23] = irqo;
  assign \apbo[prdata] [22] = irqo;
  assign \apbo[prdata] [21] = irqo;
  assign \apbo[prdata] [20] = irqo;
  assign \apbo[prdata] [19] = irqo;
  assign \apbo[prdata] [18] = irqo;
  assign \apbo[prdata] [17] = irqo;
  assign \apbo[prdata] [16] = irqo;
  assign \apbo[prdata] [15:0] = \^apbo[prdata] [15:0];
  assign \irqo[0][index] [3] = irqo;
  assign \irqo[0][index] [2] = irqo;
  assign \irqo[0][index] [1] = irqo;
  assign \irqo[0][index] [0] = irqo;
  assign \irqo[0][pwdnewaddr] [31:2] = \irqo[3][pwdnewaddr] ;
  assign \irqo[0][pwdsetaddr]  = \irqo[0][svtclrtt] ;
  assign \irqo[0][rstrun]  = \^irqo[3][index] [1];
  assign \irqo[0][rstvec] [31] = irqo;
  assign \irqo[0][rstvec] [30] = irqo;
  assign \irqo[0][rstvec] [29] = irqo;
  assign \irqo[0][rstvec] [28] = irqo;
  assign \irqo[0][rstvec] [27] = irqo;
  assign \irqo[0][rstvec] [26] = irqo;
  assign \irqo[0][rstvec] [25] = irqo;
  assign \irqo[0][rstvec] [24] = irqo;
  assign \irqo[0][rstvec] [23] = irqo;
  assign \irqo[0][rstvec] [22] = irqo;
  assign \irqo[0][rstvec] [21] = irqo;
  assign \irqo[0][rstvec] [20] = irqo;
  assign \irqo[0][rstvec] [19] = irqo;
  assign \irqo[0][rstvec] [18] = irqo;
  assign \irqo[0][rstvec] [17] = irqo;
  assign \irqo[0][rstvec] [16] = irqo;
  assign \irqo[0][rstvec] [15] = irqo;
  assign \irqo[0][rstvec] [14] = irqo;
  assign \irqo[0][rstvec] [13] = irqo;
  assign \irqo[0][rstvec] [12] = irqo;
  assign \irqo[1][index] [3] = irqo;
  assign \irqo[1][index] [2] = irqo;
  assign \irqo[1][index] [1] = irqo;
  assign \irqo[1][index] [0] = \^irqo[3][index] [1];
  assign \irqo[1][pwdnewaddr] [31:2] = \irqo[3][pwdnewaddr] ;
  assign \irqo[1][pwdsetaddr]  = \irqo[1][svtclrtt] ;
  assign \irqo[1][rstrun]  = irqo;
  assign \irqo[1][rstvec] [31] = irqo;
  assign \irqo[1][rstvec] [30] = irqo;
  assign \irqo[1][rstvec] [29] = irqo;
  assign \irqo[1][rstvec] [28] = irqo;
  assign \irqo[1][rstvec] [27] = irqo;
  assign \irqo[1][rstvec] [26] = irqo;
  assign \irqo[1][rstvec] [25] = irqo;
  assign \irqo[1][rstvec] [24] = irqo;
  assign \irqo[1][rstvec] [23] = irqo;
  assign \irqo[1][rstvec] [22] = irqo;
  assign \irqo[1][rstvec] [21] = irqo;
  assign \irqo[1][rstvec] [20] = irqo;
  assign \irqo[1][rstvec] [19] = irqo;
  assign \irqo[1][rstvec] [18] = irqo;
  assign \irqo[1][rstvec] [17] = irqo;
  assign \irqo[1][rstvec] [16] = irqo;
  assign \irqo[1][rstvec] [15] = irqo;
  assign \irqo[1][rstvec] [14] = irqo;
  assign \irqo[1][rstvec] [13] = irqo;
  assign \irqo[1][rstvec] [12] = irqo;
  assign \irqo[2][index] [3] = irqo;
  assign \irqo[2][index] [2] = irqo;
  assign \irqo[2][index] [1] = \^irqo[3][index] [1];
  assign \irqo[2][index] [0] = irqo;
  assign \irqo[2][pwdnewaddr] [31:2] = \irqo[3][pwdnewaddr] ;
  assign \irqo[2][pwdsetaddr]  = \irqo[2][svtclrtt] ;
  assign \irqo[2][rstrun]  = irqo;
  assign \irqo[2][rstvec] [31] = irqo;
  assign \irqo[2][rstvec] [30] = irqo;
  assign \irqo[2][rstvec] [29] = irqo;
  assign \irqo[2][rstvec] [28] = irqo;
  assign \irqo[2][rstvec] [27] = irqo;
  assign \irqo[2][rstvec] [26] = irqo;
  assign \irqo[2][rstvec] [25] = irqo;
  assign \irqo[2][rstvec] [24] = irqo;
  assign \irqo[2][rstvec] [23] = irqo;
  assign \irqo[2][rstvec] [22] = irqo;
  assign \irqo[2][rstvec] [21] = irqo;
  assign \irqo[2][rstvec] [20] = irqo;
  assign \irqo[2][rstvec] [19] = irqo;
  assign \irqo[2][rstvec] [18] = irqo;
  assign \irqo[2][rstvec] [17] = irqo;
  assign \irqo[2][rstvec] [16] = irqo;
  assign \irqo[2][rstvec] [15] = irqo;
  assign \irqo[2][rstvec] [14] = irqo;
  assign \irqo[2][rstvec] [13] = irqo;
  assign \irqo[2][rstvec] [12] = irqo;
  assign \irqo[3][index] [3] = irqo;
  assign \irqo[3][index] [2] = irqo;
  assign \irqo[3][index] [1] = \^irqo[3][index] [1];
  assign \irqo[3][index] [0] = \^irqo[3][index] [1];
  assign \irqo[3][pwdsetaddr]  = \irqo[3][svtclrtt] ;
  assign \irqo[3][rstrun]  = irqo;
  assign \irqo[3][rstvec] [31] = irqo;
  assign \irqo[3][rstvec] [30] = irqo;
  assign \irqo[3][rstvec] [29] = irqo;
  assign \irqo[3][rstvec] [28] = irqo;
  assign \irqo[3][rstvec] [27] = irqo;
  assign \irqo[3][rstvec] [26] = irqo;
  assign \irqo[3][rstvec] [25] = irqo;
  assign \irqo[3][rstvec] [24] = irqo;
  assign \irqo[3][rstvec] [23] = irqo;
  assign \irqo[3][rstvec] [22] = irqo;
  assign \irqo[3][rstvec] [21] = irqo;
  assign \irqo[3][rstvec] [20] = irqo;
  assign \irqo[3][rstvec] [19] = irqo;
  assign \irqo[3][rstvec] [18] = irqo;
  assign \irqo[3][rstvec] [17] = irqo;
  assign \irqo[3][rstvec] [16] = irqo;
  assign \irqo[3][rstvec] [15] = irqo;
  assign \irqo[3][rstvec] [14] = irqo;
  assign \irqo[3][rstvec] [13] = irqo;
  assign \irqo[3][rstvec] [12] = irqo;
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\^irqo[3][index] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \apbo[prdata][0]_INST_0 
       (.I0(\irqi[0][pwd] ),
        .I1(\apbi[paddr] [3]),
        .I2(\irqi[0][err] ),
        .I3(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .O(\^apbo[prdata] [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFB)) 
    \apbo[prdata][0]_INST_0_i_1 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [6]),
        .I3(\apbi[paddr] [7]),
        .O(\apbo[prdata][0]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][10]_INST_0 
       (.I0(\apbo[prdata][10]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][10]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [10]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][10]_INST_0_i_1 
       (.I0(\apbo[prdata][10]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in14_in),
        .I4(\apbo[prdata][10]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][10]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][10]_INST_0_i_2 
       (.I0(\apbo[prdata][10]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [9]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [9]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][10]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][10]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [9]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [9]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][10]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][10]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][10]_INST_0_i_4 
       (.I0(p_6_in[10]),
        .I1(p_5_in[10]),
        .I2(\r_reg[iforce][0]__0 [9]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][10]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][10]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [9]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [9]),
        .O(\apbo[prdata][10]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][10]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [9]),
        .I1(\r_reg[iforce][0]__0 [9]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][10]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][11]_INST_0 
       (.I0(\apbo[prdata][11]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][11]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [11]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][11]_INST_0_i_1 
       (.I0(\apbo[prdata][11]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in12_in),
        .I4(\apbo[prdata][11]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][11]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][11]_INST_0_i_2 
       (.I0(\apbo[prdata][11]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [10]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [10]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][11]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][11]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [10]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [10]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][11]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][11]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][11]_INST_0_i_4 
       (.I0(p_6_in[11]),
        .I1(p_5_in[11]),
        .I2(\r_reg[iforce][0]__0 [10]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][11]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][11]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [10]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [10]),
        .O(\apbo[prdata][11]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][11]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [10]),
        .I1(\r_reg[iforce][0]__0 [10]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][11]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][12]_INST_0 
       (.I0(\apbo[prdata][12]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][12]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [12]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][12]_INST_0_i_1 
       (.I0(\apbo[prdata][12]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in10_in),
        .I4(\apbo[prdata][12]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][12]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][12]_INST_0_i_2 
       (.I0(\apbo[prdata][12]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [11]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [11]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][12]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][12]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [11]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [11]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][12]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][12]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][12]_INST_0_i_4 
       (.I0(p_6_in[12]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][0]__0 [11]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][12]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][12]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [11]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [11]),
        .O(\apbo[prdata][12]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][12]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [11]),
        .I1(\r_reg[iforce][0]__0 [11]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][12]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][13]_INST_0 
       (.I0(\apbo[prdata][13]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][13]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [13]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][13]_INST_0_i_1 
       (.I0(\apbo[prdata][13]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in8_in),
        .I4(\apbo[prdata][13]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][13]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][13]_INST_0_i_2 
       (.I0(\apbo[prdata][13]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [12]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [12]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][13]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][13]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [12]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [12]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][13]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][13]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][13]_INST_0_i_4 
       (.I0(p_6_in[13]),
        .I1(p_5_in[13]),
        .I2(\r_reg[iforce][0]__0 [12]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][13]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][13]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [12]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [12]),
        .O(\apbo[prdata][13]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][13]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [12]),
        .I1(\r_reg[iforce][0]__0 [12]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][13]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][14]_INST_0 
       (.I0(\apbo[prdata][14]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][14]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [14]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][14]_INST_0_i_1 
       (.I0(\apbo[prdata][14]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in6_in),
        .I4(\apbo[prdata][14]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][14]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][14]_INST_0_i_2 
       (.I0(\apbo[prdata][14]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [13]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [13]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][14]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][14]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [13]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [13]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][14]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][14]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][14]_INST_0_i_4 
       (.I0(p_6_in[14]),
        .I1(p_5_in[14]),
        .I2(\r_reg[iforce][0]__0 [13]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][14]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][14]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [13]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [13]),
        .O(\apbo[prdata][14]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][14]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [13]),
        .I1(\r_reg[iforce][0]__0 [13]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][14]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][15]_INST_0 
       (.I0(\apbo[prdata][15]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [15]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][15]_INST_0_i_1 
       (.I0(\apbo[prdata][15]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in4_in),
        .I4(\apbo[prdata][15]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata][15]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][15]_INST_0_i_2 
       (.I0(\apbo[prdata][15]_INST_0_i_6_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [14]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [14]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][15]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][15]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [14]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [14]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][15]_INST_0_i_8_n_0 ),
        .O(\apbo[prdata][15]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \apbo[prdata][15]_INST_0_i_4 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [4]),
        .O(\apbo[prdata][15]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][15]_INST_0_i_5 
       (.I0(p_6_in[15]),
        .I1(p_5_in[15]),
        .I2(\r_reg[iforce][0]__0 [14]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][15]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][15]_INST_0_i_6 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [14]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [14]),
        .O(\apbo[prdata][15]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \apbo[prdata][15]_INST_0_i_7 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [4]),
        .O(\apbo[prdata][15]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][15]_INST_0_i_8 
       (.I0(\r_reg[iforce][2]__0 [14]),
        .I1(\r_reg[iforce][0]__0 [14]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][15]_INST_0_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \apbo[prdata][1]_INST_0 
       (.I0(\apbo[prdata][1]_INST_0_i_1_n_0 ),
        .I1(\apbi[paddr] [6]),
        .I2(\apbo[prdata][1]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbo[prdata][1]_INST_0_i_3_n_0 ),
        .O(\^apbo[prdata] [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][1]_INST_0_i_1 
       (.I0(\apbo[prdata][1]_INST_0_i_4_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [0]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [0]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][1]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][1]_INST_0_i_2 
       (.I0(\r_reg[iforce][3]__0 [0]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [0]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][1]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata][1]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F33BFB30C008C80)) 
    \apbo[prdata][1]_INST_0_i_3 
       (.I0(\irqi[1][err] ),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbo[prdata][1]_INST_0_i_6_n_0 ),
        .I4(\apbi[paddr] [2]),
        .I5(\apbo[prdata][1]_INST_0_i_7_n_0 ),
        .O(\apbo[prdata][1]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][1]_INST_0_i_4 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [0]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [0]),
        .O(\apbo[prdata][1]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][1]_INST_0_i_5 
       (.I0(\r_reg[iforce][2]__0 [0]),
        .I1(\r_reg[iforce][0]__0 [0]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][1]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF2000)) 
    \apbo[prdata][1]_INST_0_i_6 
       (.I0(\r_reg[ibroadcast_n_0_][1] ),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [4]),
        .I4(\irqi[1][pwd] ),
        .O(\apbo[prdata][1]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \apbo[prdata][1]_INST_0_i_7 
       (.I0(\r_reg[iforce][0]__0 [0]),
        .I1(\apbi[paddr] [3]),
        .I2(p_5_in[1]),
        .I3(\apbi[paddr] [2]),
        .I4(p_6_in[1]),
        .O(\apbo[prdata][1]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \apbo[prdata][26]_INST_0 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [6]),
        .I3(\apbi[paddr] [7]),
        .O(\^apbo[prdata] [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \apbo[prdata][27]_INST_0 
       (.I0(\apbi[paddr] [7]),
        .I1(\apbi[paddr] [6]),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [2]),
        .O(apbo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \apbo[prdata][2]_INST_0 
       (.I0(\apbo[prdata][2]_INST_0_i_1_n_0 ),
        .I1(\apbi[paddr] [6]),
        .I2(\apbo[prdata][2]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbo[prdata][2]_INST_0_i_3_n_0 ),
        .O(\^apbo[prdata] [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][2]_INST_0_i_1 
       (.I0(\apbo[prdata][2]_INST_0_i_4_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [1]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [1]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][2]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][2]_INST_0_i_2 
       (.I0(\r_reg[iforce][3]__0 [1]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [1]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][2]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata][2]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F33BFB30C008C80)) 
    \apbo[prdata][2]_INST_0_i_3 
       (.I0(\irqi[2][err] ),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbo[prdata][2]_INST_0_i_6_n_0 ),
        .I4(\apbi[paddr] [2]),
        .I5(\apbo[prdata][2]_INST_0_i_7_n_0 ),
        .O(\apbo[prdata][2]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][2]_INST_0_i_4 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [1]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [1]),
        .O(\apbo[prdata][2]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][2]_INST_0_i_5 
       (.I0(\r_reg[iforce][2]__0 [1]),
        .I1(\r_reg[iforce][0]__0 [1]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][2]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF2000)) 
    \apbo[prdata][2]_INST_0_i_6 
       (.I0(p_0_in30_in),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [4]),
        .I4(\irqi[2][pwd] ),
        .O(\apbo[prdata][2]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \apbo[prdata][2]_INST_0_i_7 
       (.I0(\r_reg[iforce][0]__0 [1]),
        .I1(\apbi[paddr] [3]),
        .I2(p_5_in[2]),
        .I3(\apbi[paddr] [2]),
        .I4(p_6_in[2]),
        .O(\apbo[prdata][2]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \apbo[prdata][3]_INST_0 
       (.I0(\apbo[prdata][3]_INST_0_i_1_n_0 ),
        .I1(\apbi[paddr] [6]),
        .I2(\apbo[prdata][3]_INST_0_i_2_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbo[prdata][3]_INST_0_i_3_n_0 ),
        .O(\^apbo[prdata] [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][3]_INST_0_i_1 
       (.I0(\apbo[prdata][3]_INST_0_i_4_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [2]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][3]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][3]_INST_0_i_2 
       (.I0(\r_reg[iforce][3]__0 [2]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [2]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][3]_INST_0_i_5_n_0 ),
        .O(\apbo[prdata][3]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3F33BFB30C008C80)) 
    \apbo[prdata][3]_INST_0_i_3 
       (.I0(\irqi[3][err] ),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbo[prdata][3]_INST_0_i_6_n_0 ),
        .I4(\apbi[paddr] [2]),
        .I5(\apbo[prdata][3]_INST_0_i_7_n_0 ),
        .O(\apbo[prdata][3]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][3]_INST_0_i_4 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [2]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [2]),
        .O(\apbo[prdata][3]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][3]_INST_0_i_5 
       (.I0(\r_reg[iforce][2]__0 [2]),
        .I1(\r_reg[iforce][0]__0 [2]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][3]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF2000)) 
    \apbo[prdata][3]_INST_0_i_6 
       (.I0(p_0_in28_in),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [4]),
        .I4(\irqi[3][pwd] ),
        .O(\apbo[prdata][3]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \apbo[prdata][3]_INST_0_i_7 
       (.I0(\r_reg[iforce][0]__0 [2]),
        .I1(\apbi[paddr] [3]),
        .I2(p_5_in[3]),
        .I3(\apbi[paddr] [2]),
        .I4(p_6_in[3]),
        .O(\apbo[prdata][3]_INST_0_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][4]_INST_0 
       (.I0(\apbo[prdata][4]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][4]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [4]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][4]_INST_0_i_1 
       (.I0(\apbo[prdata][4]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in26_in),
        .I4(\apbo[prdata][4]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][4]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][4]_INST_0_i_2 
       (.I0(\apbo[prdata][4]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [3]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [3]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][4]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][4]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [3]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [3]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][4]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][4]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][4]_INST_0_i_4 
       (.I0(p_6_in[4]),
        .I1(p_5_in[4]),
        .I2(\r_reg[iforce][0]__0 [3]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][4]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][4]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [3]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [3]),
        .O(\apbo[prdata][4]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][4]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [3]),
        .I1(\r_reg[iforce][0]__0 [3]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][4]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][5]_INST_0 
       (.I0(\apbo[prdata][5]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][5]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [5]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][5]_INST_0_i_1 
       (.I0(\apbo[prdata][5]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in24_in),
        .I4(\apbo[prdata][5]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][5]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][5]_INST_0_i_2 
       (.I0(\apbo[prdata][5]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [4]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [4]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][5]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][5]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [4]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [4]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][5]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][5]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][5]_INST_0_i_4 
       (.I0(p_6_in[5]),
        .I1(p_5_in[5]),
        .I2(\r_reg[iforce][0]__0 [4]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][5]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][5]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [4]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [4]),
        .O(\apbo[prdata][5]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][5]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [4]),
        .I1(\r_reg[iforce][0]__0 [4]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][5]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][6]_INST_0 
       (.I0(\apbo[prdata][6]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][6]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [6]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][6]_INST_0_i_1 
       (.I0(\apbo[prdata][6]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in22_in),
        .I4(\apbo[prdata][6]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][6]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][6]_INST_0_i_2 
       (.I0(\apbo[prdata][6]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [5]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][6]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][6]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [5]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [5]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][6]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][6]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][6]_INST_0_i_4 
       (.I0(p_6_in[6]),
        .I1(p_5_in[6]),
        .I2(\r_reg[iforce][0]__0 [5]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][6]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][6]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [5]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [5]),
        .O(\apbo[prdata][6]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][6]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [5]),
        .I1(\r_reg[iforce][0]__0 [5]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][6]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][7]_INST_0 
       (.I0(\apbo[prdata][7]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][7]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [7]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][7]_INST_0_i_1 
       (.I0(\apbo[prdata][7]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in20_in),
        .I4(\apbo[prdata][7]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][7]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][7]_INST_0_i_2 
       (.I0(\apbo[prdata][7]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [6]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [6]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][7]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][7]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [6]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [6]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][7]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][7]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][7]_INST_0_i_4 
       (.I0(p_6_in[7]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][0]__0 [6]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][7]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][7]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [6]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [6]),
        .O(\apbo[prdata][7]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][7]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [6]),
        .I1(\r_reg[iforce][0]__0 [6]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][7]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][8]_INST_0 
       (.I0(\apbo[prdata][8]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][8]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [8]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][8]_INST_0_i_1 
       (.I0(\apbo[prdata][8]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in18_in),
        .I4(\apbo[prdata][8]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][8]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][8]_INST_0_i_2 
       (.I0(\apbo[prdata][8]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [7]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [7]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][8]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][8]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [7]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [7]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][8]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][8]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][8]_INST_0_i_4 
       (.I0(p_6_in[8]),
        .I1(p_5_in[8]),
        .I2(\r_reg[iforce][0]__0 [7]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][8]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][8]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [7]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [7]),
        .O(\apbo[prdata][8]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][8]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [7]),
        .I1(\r_reg[iforce][0]__0 [7]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][8]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \apbo[prdata][9]_INST_0 
       (.I0(\apbo[prdata][9]_INST_0_i_1_n_0 ),
        .I1(\apbo[prdata][9]_INST_0_i_2_n_0 ),
        .O(\^apbo[prdata] [9]),
        .S(\apbi[paddr] [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBBBBB888)) 
    \apbo[prdata][9]_INST_0_i_1 
       (.I0(\apbo[prdata][9]_INST_0_i_3_n_0 ),
        .I1(\apbi[paddr] [7]),
        .I2(\apbo[prdata][15]_INST_0_i_4_n_0 ),
        .I3(p_0_in16_in),
        .I4(\apbo[prdata][9]_INST_0_i_4_n_0 ),
        .O(\apbo[prdata][9]_INST_0_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE222E2)) 
    \apbo[prdata][9]_INST_0_i_2 
       (.I0(\apbo[prdata][9]_INST_0_i_5_n_0 ),
        .I1(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I2(\r_reg[imask][1]__0 [8]),
        .I3(\apbi[paddr] [3]),
        .I4(\r_reg[imask][3]__0 [8]),
        .I5(\apbi[paddr] [7]),
        .O(\apbo[prdata][9]_INST_0_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \apbo[prdata][9]_INST_0_i_3 
       (.I0(\r_reg[iforce][3]__0 [8]),
        .I1(\apbi[paddr] [3]),
        .I2(\r_reg[iforce][1]__0 [8]),
        .I3(\apbo[prdata][15]_INST_0_i_7_n_0 ),
        .I4(\apbo[prdata][9]_INST_0_i_6_n_0 ),
        .O(\apbo[prdata][9]_INST_0_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000F0CCAA)) 
    \apbo[prdata][9]_INST_0_i_4 
       (.I0(p_6_in[9]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][0]__0 [8]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\apbo[prdata][9]_INST_0_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000F0400000004)) 
    \apbo[prdata][9]_INST_0_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\r_reg[imask][0]__0 [8]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r_reg[imask][2]__0 [8]),
        .O(\apbo[prdata][9]_INST_0_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000000000AA0C)) 
    \apbo[prdata][9]_INST_0_i_6 
       (.I0(\r_reg[iforce][2]__0 [8]),
        .I1(\r_reg[iforce][0]__0 [8]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [5]),
        .O(\apbo[prdata][9]_INST_0_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'hFFFFFF0E)) 
    \r[clkcount][0]_i_1 
       (.I0(\r_reg[clkcount_n_0_][2] ),
        .I1(\r_reg[clkcount_n_0_][1] ),
        .I2(r_reg),
        .I3(\r[clkcount][2]_i_2_n_0 ),
        .I4(v),
        .O(r));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFC2)) 
    \r[clkcount][1]_i_1 
       (.I0(\r_reg[clkcount_n_0_][2] ),
        .I1(\r_reg[clkcount_n_0_][1] ),
        .I2(r_reg),
        .I3(\r[clkcount][2]_i_2_n_0 ),
        .I4(v),
        .O(\r[clkcount][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'hFFFFFFA8)) 
    \r[clkcount][2]_i_1 
       (.I0(\r_reg[clkcount_n_0_][2] ),
        .I1(\r_reg[clkcount_n_0_][1] ),
        .I2(r_reg),
        .I3(\r[clkcount][2]_i_2_n_0 ),
        .I4(v),
        .O(\r[clkcount][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000008)) 
    \r[clkcount][2]_i_2 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\r[cpurst][0]_i_3_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [2]),
        .I5(\apbi[paddr] [6]),
        .O(\r[clkcount][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444444444F44)) 
    \r[cpurst][0]_i_1 
       (.I0(\r[cpurst][0]_i_2_n_0 ),
        .I1(\irqo[0][svtclrtt] ),
        .I2(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I3(\apbi[pwdata] [0]),
        .I4(\apbi[paddr] [3]),
        .I5(\r[cpurst][0]_i_3_n_0 ),
        .O(\v[cpurst]1_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFDFFFF)) 
    \r[cpurst][0]_i_2 
       (.I0(\irqo[3][pwdnewaddr] [2]),
        .I1(\r_reg[clkcount_n_0_][2] ),
        .I2(\r_reg[clkcount_n_0_][1] ),
        .I3(r_reg),
        .I4(\r_reg[setaddrboot_n_0_] ),
        .O(\r[cpurst][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r[cpurst][0]_i_3 
       (.I0(\apbi[penable] ),
        .I1(apbi[2]),
        .I2(\apbi[pwrite] ),
        .O(\r[cpurst][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[cpurst][1]_i_1 
       (.I0(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I1(\apbi[pwdata] [1]),
        .I2(\apbi[paddr] [3]),
        .I3(\r[cpurst][0]_i_3_n_0 ),
        .I4(\r[cpurst][0]_i_2_n_0 ),
        .I5(\irqo[1][svtclrtt] ),
        .O(\v[cpurst]1_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[cpurst][2]_i_1 
       (.I0(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I1(\apbi[pwdata] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\r[cpurst][0]_i_3_n_0 ),
        .I4(\r[cpurst][0]_i_2_n_0 ),
        .I5(\irqo[2][svtclrtt] ),
        .O(\v[cpurst]1_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100010)) 
    \r[cpurst][3]_i_1 
       (.I0(\apbi[paddr] [3]),
        .I1(\r[cpurst][0]_i_3_n_0 ),
        .I2(\apbi[pwdata] [3]),
        .I3(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I4(\r[cpurst][0]_i_2_n_0 ),
        .I5(\irqo[3][svtclrtt] ),
        .O(\v[cpurst]1_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0D0DDD0D0D0D0D0)) 
    \r[forceerr][0]_i_1 
       (.I0(\irqi[0][err] ),
        .I1(\r[forceerr][0]_i_2_n_0 ),
        .I2(\irqo[0][forceerr] ),
        .I3(\apbi[pwdata] [0]),
        .I4(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I5(\r[forceerr][0]_i_3_n_0 ),
        .O(\r[forceerr][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r[forceerr][0]_i_2 
       (.I0(\r_reg[clkcount_n_0_][2] ),
        .I1(\r_reg[clkcount_n_0_][1] ),
        .I2(r_reg),
        .O(\r[forceerr][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \r[forceerr][0]_i_3 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[pwrite] ),
        .I2(apbi[2]),
        .I3(\apbi[penable] ),
        .O(\r[forceerr][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0D0DDD0D0D0D0D0)) 
    \r[forceerr][1]_i_1 
       (.I0(\irqi[1][err] ),
        .I1(\r[forceerr][0]_i_2_n_0 ),
        .I2(\irqo[1][forceerr] ),
        .I3(\apbi[pwdata] [1]),
        .I4(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I5(\r[forceerr][0]_i_3_n_0 ),
        .O(\r[forceerr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0D0DDD0D0D0D0D0)) 
    \r[forceerr][2]_i_1 
       (.I0(\irqi[2][err] ),
        .I1(\r[forceerr][0]_i_2_n_0 ),
        .I2(\irqo[2][forceerr] ),
        .I3(\apbi[pwdata] [2]),
        .I4(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I5(\r[forceerr][0]_i_3_n_0 ),
        .O(\r[forceerr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0D0DDD0D0D0D0D0)) 
    \r[forceerr][3]_i_1 
       (.I0(\irqi[3][err] ),
        .I1(\r[forceerr][0]_i_2_n_0 ),
        .I2(\irqo[3][forceerr] ),
        .I3(\r[forceerr][0]_i_3_n_0 ),
        .I4(\apbo[prdata][0]_INST_0_i_1_n_0 ),
        .I5(\apbi[pwdata] [3]),
        .O(\r[forceerr][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001000000000)) 
    \r[ibroadcast][15]_i_1 
       (.I0(\apbi[paddr] [7]),
        .I1(\apbi[paddr] [6]),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [3]),
        .I4(\r[cpurst][0]_i_3_n_0 ),
        .I5(\apbi[paddr] [2]),
        .O(\v[ibroadcast] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFBFFFFF)) 
    \r[iforce][0][10]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][10]_i_2_n_0 ),
        .O(\r[iforce][0][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][10]_i_2 
       (.I0(\r_reg[iforce][0]__0 [9]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [26]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][10]_i_3_n_0 ),
        .O(\r[iforce][0][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][10]_i_3 
       (.I0(\r[iforce][3][10]_i_2_n_0 ),
        .I1(\apbi[pwdata] [10]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [26]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BFFFFFFF)) 
    \r[iforce][0][11]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][11]_i_2_n_0 ),
        .O(\r[iforce][0][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][11]_i_2 
       (.I0(\r_reg[iforce][0]__0 [10]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [27]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][11]_i_3_n_0 ),
        .O(\r[iforce][0][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][11]_i_3 
       (.I0(\r[iforce][3][11]_i_2_n_0 ),
        .I1(\apbi[pwdata] [11]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [27]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EFFFFFFF)) 
    \r[iforce][0][12]_i_1 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(irqi),
        .I3(\irqi[0][irl] [3]),
        .I4(\irqi[0][irl] [2]),
        .I5(\r[iforce][0][12]_i_2_n_0 ),
        .O(\r[iforce][0][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][12]_i_2 
       (.I0(\r_reg[iforce][0]__0 [11]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [28]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][12]_i_3_n_0 ),
        .O(\r[iforce][0][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][12]_i_3 
       (.I0(\r[iforce][3][12]_i_2_n_0 ),
        .I1(\apbi[pwdata] [12]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [28]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BFFFFFFF)) 
    \r[iforce][0][13]_i_1 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(irqi),
        .I3(\irqi[0][irl] [3]),
        .I4(\irqi[0][irl] [2]),
        .I5(\r[iforce][0][13]_i_2_n_0 ),
        .O(\r[iforce][0][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][13]_i_2 
       (.I0(\r_reg[iforce][0]__0 [12]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [29]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][13]_i_3_n_0 ),
        .O(\r[iforce][0][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][13]_i_3 
       (.I0(\r[iforce][3][13]_i_2_n_0 ),
        .I1(\apbi[pwdata] [13]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [29]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BFFFFFFF)) 
    \r[iforce][0][14]_i_1 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(irqi),
        .I3(\irqi[0][irl] [3]),
        .I4(\irqi[0][irl] [2]),
        .I5(\r[iforce][0][14]_i_2_n_0 ),
        .O(\r[iforce][0][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][14]_i_2 
       (.I0(\r_reg[iforce][0]__0 [13]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [30]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][14]_i_3_n_0 ),
        .O(\r[iforce][0][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00088888)) 
    \r[iforce][0][14]_i_3 
       (.I0(\apbi[pwdata] [14]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\r[iforce][0][15]_i_4_n_0 ),
        .I3(\apbi[pwdata] [30]),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][3][14]_i_3_n_0 ),
        .O(\r[iforce][0][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000007FFFFFFF)) 
    \r[iforce][0][15]_i_1 
       (.I0(irqi),
        .I1(\irqi[0][irl] [3]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][15]_i_2_n_0 ),
        .O(\r[iforce][0][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][15]_i_2 
       (.I0(\r_reg[iforce][0]__0 [14]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [31]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][15]_i_5_n_0 ),
        .O(\r[iforce][0][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1111111100000100)) 
    \r[iforce][0][15]_i_3 
       (.I0(\r[cpurst][0]_i_3_n_0 ),
        .I1(\apbi[paddr] [6]),
        .I2(\apbi[paddr] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[iforce][0][15]_i_4 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [5]),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [3]),
        .O(\r[iforce][0][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00088888)) 
    \r[iforce][0][15]_i_5 
       (.I0(\apbi[pwdata] [15]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\r[iforce][0][15]_i_4_n_0 ),
        .I3(\apbi[pwdata] [31]),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][1][15]_i_3_n_0 ),
        .O(\r[iforce][0][15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFBFFFF)) 
    \r[iforce][0][1]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .I5(\r[iforce][0][1]_i_2_n_0 ),
        .O(\r[iforce][0][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][1]_i_2 
       (.I0(\r_reg[iforce][0]__0 [0]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [17]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][1]_i_3_n_0 ),
        .O(\r[iforce][0][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][1]_i_3 
       (.I0(\r[iforce][3][1]_i_2_n_0 ),
        .I1(\apbi[pwdata] [1]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [17]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFBFFFF)) 
    \r[iforce][0][2]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][2]_i_2_n_0 ),
        .O(\r[iforce][0][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][2]_i_2 
       (.I0(\r_reg[iforce][0]__0 [1]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [18]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][2]_i_3_n_0 ),
        .O(\r[iforce][0][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][2]_i_3 
       (.I0(\r[iforce][3][2]_i_2_n_0 ),
        .I1(\apbi[pwdata] [2]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [18]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FBFFFFFF)) 
    \r[iforce][0][3]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][3]_i_2_n_0 ),
        .O(\r[iforce][0][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][3]_i_2 
       (.I0(\r_reg[iforce][0]__0 [2]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [19]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][3]_i_3_n_0 ),
        .O(\r[iforce][0][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][3]_i_3 
       (.I0(\r[iforce][3][3]_i_2_n_0 ),
        .I1(\apbi[pwdata] [3]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [19]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFEFFFFF)) 
    \r[iforce][0][4]_i_1 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(irqi),
        .I3(\irqi[0][irl] [3]),
        .I4(\irqi[0][irl] [2]),
        .I5(\r[iforce][0][4]_i_2_n_0 ),
        .O(\r[iforce][0][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][4]_i_2 
       (.I0(\r_reg[iforce][0]__0 [3]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [20]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][4]_i_3_n_0 ),
        .O(\r[iforce][0][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][4]_i_3 
       (.I0(\r[iforce][3][4]_i_2_n_0 ),
        .I1(\apbi[pwdata] [4]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [20]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFDFFFFF)) 
    \r[iforce][0][5]_i_1 
       (.I0(irqi),
        .I1(\irqi[0][irl] [3]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .I5(\r[iforce][0][5]_i_2_n_0 ),
        .O(\r[iforce][0][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][5]_i_2 
       (.I0(\r_reg[iforce][0]__0 [4]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [21]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][5]_i_3_n_0 ),
        .O(\r[iforce][0][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][5]_i_3 
       (.I0(\r[iforce][3][5]_i_2_n_0 ),
        .I1(\apbi[pwdata] [5]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [21]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFDFFFFF)) 
    \r[iforce][0][6]_i_1 
       (.I0(irqi),
        .I1(\irqi[0][irl] [3]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][6]_i_2_n_0 ),
        .O(\r[iforce][0][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][6]_i_2 
       (.I0(\r_reg[iforce][0]__0 [5]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [22]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][6]_i_3_n_0 ),
        .O(\r[iforce][0][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][6]_i_3 
       (.I0(\r[iforce][3][6]_i_2_n_0 ),
        .I1(\apbi[pwdata] [6]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [22]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000DFFFFFFF)) 
    \r[iforce][0][7]_i_1 
       (.I0(irqi),
        .I1(\irqi[0][irl] [3]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .I5(\r[iforce][0][7]_i_2_n_0 ),
        .O(\r[iforce][0][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][7]_i_2 
       (.I0(\r_reg[iforce][0]__0 [6]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [23]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][7]_i_3_n_0 ),
        .O(\r[iforce][0][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][7]_i_3 
       (.I0(\r[iforce][3][7]_i_2_n_0 ),
        .I1(\apbi[pwdata] [7]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [23]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAA8AAA)) 
    \r[iforce][0][8]_i_1 
       (.I0(\r[iforce][0][8]_i_2_n_0 ),
        .I1(\irqi[0][irl] [2]),
        .I2(irqi),
        .I3(\irqi[0][irl] [3]),
        .I4(\irqi[0][irl] [0]),
        .I5(\irqi[0][irl] [1]),
        .O(\r[iforce][0][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFF7550000)) 
    \r[iforce][0][8]_i_2 
       (.I0(\r[iforce][0][15]_i_3_n_0 ),
        .I1(\apbi[pwdata] [24]),
        .I2(\r[iforce][0][15]_i_4_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\r_reg[iforce][0]__0 [7]),
        .I5(\r[iforce][0][8]_i_3_n_0 ),
        .O(\r[iforce][0][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][8]_i_3 
       (.I0(\r[iforce][3][8]_i_2_n_0 ),
        .I1(\apbi[pwdata] [8]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [24]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFBFFFFF)) 
    \r[iforce][0][9]_i_1 
       (.I0(\irqi[0][irl] [2]),
        .I1(irqi),
        .I2(\irqi[0][irl] [3]),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .I5(\r[iforce][0][9]_i_2_n_0 ),
        .O(\r[iforce][0][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000055D5DDDD)) 
    \r[iforce][0][9]_i_2 
       (.I0(\r_reg[iforce][0]__0 [8]),
        .I1(\r[iforce][0][15]_i_3_n_0 ),
        .I2(\apbi[pwdata] [25]),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[paddr] [7]),
        .I5(\r[iforce][0][9]_i_3_n_0 ),
        .O(\r[iforce][0][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAEAEAEAEAEA)) 
    \r[iforce][0][9]_i_3 
       (.I0(\r[iforce][3][9]_i_2_n_0 ),
        .I1(\apbi[pwdata] [9]),
        .I2(\r[iforce][0][15]_i_3_n_0 ),
        .I3(\r[iforce][0][15]_i_4_n_0 ),
        .I4(\apbi[pwdata] [25]),
        .I5(\apbi[paddr] [7]),
        .O(\r[iforce][0][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][10]_i_1 
       (.I0(\apbi[pwdata] [10]),
        .I1(\r_reg[iforce][1]__0 [9]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [26]),
        .I4(\r[iforce][3][10]_i_2_n_0 ),
        .I5(\r[iforce][1][10]_i_2_n_0 ),
        .O(\r[iforce][1][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][1][10]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][11]_i_1 
       (.I0(\apbi[pwdata] [11]),
        .I1(\r_reg[iforce][1]__0 [10]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [27]),
        .I4(\r[iforce][3][11]_i_2_n_0 ),
        .I5(\r[iforce][1][11]_i_2_n_0 ),
        .O(\r[iforce][1][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][1][11]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][12]_i_1 
       (.I0(\apbi[pwdata] [12]),
        .I1(\r_reg[iforce][1]__0 [11]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [28]),
        .I4(\r[iforce][3][12]_i_2_n_0 ),
        .I5(\r[iforce][1][12]_i_2_n_0 ),
        .O(\r[iforce][1][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \r[iforce][1][12]_i_2 
       (.I0(\irqi[1][irl] [2]),
        .I1(\irqi[1][irl] [3]),
        .I2(\irqi[1][intack] ),
        .I3(\irqi[1][irl] [1]),
        .I4(\irqi[1][irl] [0]),
        .O(\r[iforce][1][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][13]_i_1 
       (.I0(\apbi[pwdata] [13]),
        .I1(\r_reg[iforce][1]__0 [12]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [29]),
        .I4(\r[iforce][3][13]_i_2_n_0 ),
        .I5(\r[iforce][1][13]_i_2_n_0 ),
        .O(\r[iforce][1][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][1][13]_i_2 
       (.I0(\irqi[1][irl] [2]),
        .I1(\irqi[1][irl] [3]),
        .I2(\irqi[1][intack] ),
        .I3(\irqi[1][irl] [0]),
        .I4(\irqi[1][irl] [1]),
        .O(\r[iforce][1][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][14]_i_1 
       (.I0(\apbi[pwdata] [14]),
        .I1(\r_reg[iforce][1]__0 [13]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [30]),
        .I4(\r[iforce][3][14]_i_3_n_0 ),
        .I5(\r[iforce][1][14]_i_2_n_0 ),
        .O(\r[iforce][1][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][1][14]_i_2 
       (.I0(\irqi[1][irl] [2]),
        .I1(\irqi[1][irl] [3]),
        .I2(\irqi[1][intack] ),
        .I3(\irqi[1][irl] [1]),
        .I4(\irqi[1][irl] [0]),
        .O(\r[iforce][1][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][15]_i_1 
       (.I0(\apbi[pwdata] [15]),
        .I1(\r_reg[iforce][1]__0 [14]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [31]),
        .I4(\r[iforce][1][15]_i_3_n_0 ),
        .I5(\r[iforce][1][15]_i_4_n_0 ),
        .O(\r[iforce][1][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEF)) 
    \r[iforce][1][15]_i_2 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\r[iforce][3][15]_i_4_n_0 ),
        .O(\r[iforce][1][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][1][15]_i_3 
       (.I0(\apbi[pirq] [15]),
        .I1(p_0_in4_in),
        .O(\r[iforce][1][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[iforce][1][15]_i_4 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [2]),
        .I3(\irqi[1][irl] [3]),
        .I4(\irqi[1][intack] ),
        .O(\r[iforce][1][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][1]_i_1 
       (.I0(\apbi[pwdata] [1]),
        .I1(\r_reg[iforce][1]__0 [0]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [17]),
        .I4(\r[iforce][3][1]_i_2_n_0 ),
        .I5(\r[iforce][1][1]_i_2_n_0 ),
        .O(\r[iforce][1][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][1][1]_i_2 
       (.I0(\irqi[1][irl] [0]),
        .I1(\irqi[1][irl] [1]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][2]_i_1 
       (.I0(\apbi[pwdata] [2]),
        .I1(\r_reg[iforce][1]__0 [1]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [18]),
        .I4(\r[iforce][3][2]_i_2_n_0 ),
        .I5(\r[iforce][1][2]_i_2_n_0 ),
        .O(\r[iforce][1][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][1][2]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][3]_i_1 
       (.I0(\apbi[pwdata] [3]),
        .I1(\r_reg[iforce][1]__0 [2]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [19]),
        .I4(\r[iforce][3][3]_i_2_n_0 ),
        .I5(\r[iforce][1][3]_i_2_n_0 ),
        .O(\r[iforce][1][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000800)) 
    \r[iforce][1][3]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][4]_i_1 
       (.I0(\apbi[pwdata] [4]),
        .I1(\r_reg[iforce][1]__0 [3]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [20]),
        .I4(\r[iforce][3][4]_i_2_n_0 ),
        .I5(\r[iforce][1][4]_i_2_n_0 ),
        .O(\r[iforce][1][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \r[iforce][1][4]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [2]),
        .I3(\irqi[1][irl] [3]),
        .I4(\irqi[1][intack] ),
        .O(\r[iforce][1][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][5]_i_1 
       (.I0(\apbi[pwdata] [5]),
        .I1(\r_reg[iforce][1]__0 [4]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [21]),
        .I4(\r[iforce][3][5]_i_2_n_0 ),
        .I5(\r[iforce][1][5]_i_2_n_0 ),
        .O(\r[iforce][1][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][1][5]_i_2 
       (.I0(\irqi[1][irl] [0]),
        .I1(\irqi[1][irl] [1]),
        .I2(\irqi[1][irl] [2]),
        .I3(\irqi[1][irl] [3]),
        .I4(\irqi[1][intack] ),
        .O(\r[iforce][1][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][6]_i_1 
       (.I0(\apbi[pwdata] [6]),
        .I1(\r_reg[iforce][1]__0 [5]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [22]),
        .I4(\r[iforce][3][6]_i_2_n_0 ),
        .I5(\r[iforce][1][6]_i_2_n_0 ),
        .O(\r[iforce][1][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][1][6]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [2]),
        .I3(\irqi[1][irl] [3]),
        .I4(\irqi[1][intack] ),
        .O(\r[iforce][1][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][7]_i_1 
       (.I0(\apbi[pwdata] [7]),
        .I1(\r_reg[iforce][1]__0 [6]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [23]),
        .I4(\r[iforce][3][7]_i_2_n_0 ),
        .I5(\r[iforce][1][7]_i_2_n_0 ),
        .O(\r[iforce][1][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00800000)) 
    \r[iforce][1][7]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [2]),
        .I3(\irqi[1][irl] [3]),
        .I4(\irqi[1][intack] ),
        .O(\r[iforce][1][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][8]_i_1 
       (.I0(\apbi[pwdata] [8]),
        .I1(\r_reg[iforce][1]__0 [7]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [24]),
        .I4(\r[iforce][3][8]_i_2_n_0 ),
        .I5(\r[iforce][1][8]_i_2_n_0 ),
        .O(\r[iforce][1][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \r[iforce][1][8]_i_2 
       (.I0(\irqi[1][irl] [1]),
        .I1(\irqi[1][irl] [0]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][1][9]_i_1 
       (.I0(\apbi[pwdata] [9]),
        .I1(\r_reg[iforce][1]__0 [8]),
        .I2(\r[iforce][1][15]_i_2_n_0 ),
        .I3(\apbi[pwdata] [25]),
        .I4(\r[iforce][3][9]_i_2_n_0 ),
        .I5(\r[iforce][1][9]_i_2_n_0 ),
        .O(\r[iforce][1][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][1][9]_i_2 
       (.I0(\irqi[1][irl] [0]),
        .I1(\irqi[1][irl] [1]),
        .I2(\irqi[1][irl] [3]),
        .I3(\irqi[1][intack] ),
        .I4(\irqi[1][irl] [2]),
        .O(\r[iforce][1][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][10]_i_1 
       (.I0(\apbi[pwdata] [10]),
        .I1(\r_reg[iforce][2]__0 [9]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [26]),
        .I4(\r[iforce][3][10]_i_2_n_0 ),
        .I5(\r[iforce][2][10]_i_2_n_0 ),
        .O(\r[iforce][2][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][2][10]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][11]_i_1 
       (.I0(\apbi[pwdata] [11]),
        .I1(\r_reg[iforce][2]__0 [10]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [27]),
        .I4(\r[iforce][3][11]_i_2_n_0 ),
        .I5(\r[iforce][2][11]_i_2_n_0 ),
        .O(\r[iforce][2][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][2][11]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][12]_i_1 
       (.I0(\apbi[pwdata] [12]),
        .I1(\r_reg[iforce][2]__0 [11]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [28]),
        .I4(\r[iforce][3][12]_i_2_n_0 ),
        .I5(\r[iforce][2][12]_i_2_n_0 ),
        .O(\r[iforce][2][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \r[iforce][2][12]_i_2 
       (.I0(\irqi[2][irl] [2]),
        .I1(\irqi[2][irl] [3]),
        .I2(\irqi[2][intack] ),
        .I3(\irqi[2][irl] [1]),
        .I4(\irqi[2][irl] [0]),
        .O(\r[iforce][2][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][13]_i_1 
       (.I0(\apbi[pwdata] [13]),
        .I1(\r_reg[iforce][2]__0 [12]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [29]),
        .I4(\r[iforce][3][13]_i_2_n_0 ),
        .I5(\r[iforce][2][13]_i_2_n_0 ),
        .O(\r[iforce][2][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][2][13]_i_2 
       (.I0(\irqi[2][irl] [2]),
        .I1(\irqi[2][irl] [3]),
        .I2(\irqi[2][intack] ),
        .I3(\irqi[2][irl] [0]),
        .I4(\irqi[2][irl] [1]),
        .O(\r[iforce][2][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][14]_i_1 
       (.I0(\apbi[pwdata] [14]),
        .I1(\r_reg[iforce][2]__0 [13]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [30]),
        .I4(\r[iforce][3][14]_i_3_n_0 ),
        .I5(\r[iforce][2][14]_i_3_n_0 ),
        .O(\r[iforce][2][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \r[iforce][2][14]_i_2 
       (.I0(\r[iforce][2][14]_i_4_n_0 ),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [2]),
        .O(\r[iforce][2][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][2][14]_i_3 
       (.I0(\irqi[2][irl] [2]),
        .I1(\irqi[2][irl] [3]),
        .I2(\irqi[2][intack] ),
        .I3(\irqi[2][irl] [1]),
        .I4(\irqi[2][irl] [0]),
        .O(\r[iforce][2][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBFFFFFFFFFFFFFF)) 
    \r[iforce][2][14]_i_4 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [7]),
        .I2(\apbi[paddr] [6]),
        .I3(\apbi[pwrite] ),
        .I4(apbi[2]),
        .I5(\apbi[penable] ),
        .O(\r[iforce][2][14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA00EAEAEAEAEAEA)) 
    \r[iforce][2][15]_i_1 
       (.I0(\r[iforce][2][15]_i_2_n_0 ),
        .I1(\apbi[pirq] [15]),
        .I2(p_0_in4_in),
        .I3(\r[iforce][2][15]_i_3_n_0 ),
        .I4(\irqi[2][irl] [0]),
        .I5(\irqi[2][irl] [1]),
        .O(\r[iforce][2][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCCCC0CECCCC)) 
    \r[iforce][2][15]_i_2 
       (.I0(\apbi[pwdata] [15]),
        .I1(\r_reg[iforce][2]__0 [14]),
        .I2(\r[iforce][2][15]_i_4_n_0 ),
        .I3(\apbi[pwdata] [31]),
        .I4(\apbi[paddr] [3]),
        .I5(\apbi[paddr] [4]),
        .O(\r[iforce][2][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r[iforce][2][15]_i_3 
       (.I0(\irqi[2][intack] ),
        .I1(\irqi[2][irl] [3]),
        .I2(\irqi[2][irl] [2]),
        .O(\r[iforce][2][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF8FFFF)) 
    \r[iforce][2][15]_i_4 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [2]),
        .I2(\r[cpurst][0]_i_3_n_0 ),
        .I3(\apbi[paddr] [6]),
        .I4(\apbi[paddr] [7]),
        .I5(\apbi[paddr] [5]),
        .O(\r[iforce][2][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][1]_i_1 
       (.I0(\apbi[pwdata] [1]),
        .I1(\r_reg[iforce][2]__0 [0]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [17]),
        .I4(\r[iforce][3][1]_i_2_n_0 ),
        .I5(\r[iforce][2][1]_i_2_n_0 ),
        .O(\r[iforce][2][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][2][1]_i_2 
       (.I0(\irqi[2][irl] [0]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][2]_i_1 
       (.I0(\apbi[pwdata] [2]),
        .I1(\r_reg[iforce][2]__0 [1]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [18]),
        .I4(\r[iforce][3][2]_i_2_n_0 ),
        .I5(\r[iforce][2][2]_i_2_n_0 ),
        .O(\r[iforce][2][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][2][2]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][3]_i_1 
       (.I0(\apbi[pwdata] [3]),
        .I1(\r_reg[iforce][2]__0 [2]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [19]),
        .I4(\r[iforce][3][3]_i_2_n_0 ),
        .I5(\r[iforce][2][3]_i_2_n_0 ),
        .O(\r[iforce][2][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000800)) 
    \r[iforce][2][3]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][4]_i_1 
       (.I0(\apbi[pwdata] [4]),
        .I1(\r_reg[iforce][2]__0 [3]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [20]),
        .I4(\r[iforce][3][4]_i_2_n_0 ),
        .I5(\r[iforce][2][4]_i_2_n_0 ),
        .O(\r[iforce][2][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \r[iforce][2][4]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [2]),
        .I3(\irqi[2][irl] [3]),
        .I4(\irqi[2][intack] ),
        .O(\r[iforce][2][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][5]_i_1 
       (.I0(\apbi[pwdata] [5]),
        .I1(\r_reg[iforce][2]__0 [4]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [21]),
        .I4(\r[iforce][3][5]_i_2_n_0 ),
        .I5(\r[iforce][2][5]_i_2_n_0 ),
        .O(\r[iforce][2][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][2][5]_i_2 
       (.I0(\irqi[2][irl] [0]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [2]),
        .I3(\irqi[2][irl] [3]),
        .I4(\irqi[2][intack] ),
        .O(\r[iforce][2][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][6]_i_1 
       (.I0(\apbi[pwdata] [6]),
        .I1(\r_reg[iforce][2]__0 [5]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [22]),
        .I4(\r[iforce][3][6]_i_2_n_0 ),
        .I5(\r[iforce][2][6]_i_2_n_0 ),
        .O(\r[iforce][2][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][2][6]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [2]),
        .I3(\irqi[2][irl] [3]),
        .I4(\irqi[2][intack] ),
        .O(\r[iforce][2][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][7]_i_1 
       (.I0(\apbi[pwdata] [7]),
        .I1(\r_reg[iforce][2]__0 [6]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [23]),
        .I4(\r[iforce][3][7]_i_2_n_0 ),
        .I5(\r[iforce][2][7]_i_2_n_0 ),
        .O(\r[iforce][2][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00800000)) 
    \r[iforce][2][7]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [2]),
        .I3(\irqi[2][irl] [3]),
        .I4(\irqi[2][intack] ),
        .O(\r[iforce][2][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][8]_i_1 
       (.I0(\apbi[pwdata] [8]),
        .I1(\r_reg[iforce][2]__0 [7]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [24]),
        .I4(\r[iforce][3][8]_i_2_n_0 ),
        .I5(\r[iforce][2][8]_i_2_n_0 ),
        .O(\r[iforce][2][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \r[iforce][2][8]_i_2 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][2][9]_i_1 
       (.I0(\apbi[pwdata] [9]),
        .I1(\r_reg[iforce][2]__0 [8]),
        .I2(\r[iforce][2][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [25]),
        .I4(\r[iforce][3][9]_i_2_n_0 ),
        .I5(\r[iforce][2][9]_i_2_n_0 ),
        .O(\r[iforce][2][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][2][9]_i_2 
       (.I0(\irqi[2][irl] [0]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [3]),
        .I3(\irqi[2][intack] ),
        .I4(\irqi[2][irl] [2]),
        .O(\r[iforce][2][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][10]_i_1 
       (.I0(\apbi[pwdata] [10]),
        .I1(\r_reg[iforce][3]__0 [9]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [26]),
        .I4(\r[iforce][3][10]_i_2_n_0 ),
        .I5(\r[iforce][3][10]_i_3_n_0 ),
        .O(\r[iforce][3][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][10]_i_2 
       (.I0(\apbi[pirq] [10]),
        .I1(p_0_in14_in),
        .O(\r[iforce][3][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][3][10]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][11]_i_1 
       (.I0(\apbi[pwdata] [11]),
        .I1(\r_reg[iforce][3]__0 [10]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [27]),
        .I4(\r[iforce][3][11]_i_2_n_0 ),
        .I5(\r[iforce][3][11]_i_3_n_0 ),
        .O(\r[iforce][3][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][11]_i_2 
       (.I0(\apbi[pirq] [11]),
        .I1(p_0_in12_in),
        .O(\r[iforce][3][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][3][11]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][12]_i_1 
       (.I0(\apbi[pwdata] [12]),
        .I1(\r_reg[iforce][3]__0 [11]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [28]),
        .I4(\r[iforce][3][12]_i_2_n_0 ),
        .I5(\r[iforce][3][12]_i_3_n_0 ),
        .O(\r[iforce][3][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][12]_i_2 
       (.I0(\apbi[pirq] [12]),
        .I1(p_0_in10_in),
        .O(\r[iforce][3][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \r[iforce][3][12]_i_3 
       (.I0(\irqi[3][irl] [2]),
        .I1(\irqi[3][irl] [3]),
        .I2(\irqi[3][intack] ),
        .I3(\irqi[3][irl] [1]),
        .I4(\irqi[3][irl] [0]),
        .O(\r[iforce][3][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][13]_i_1 
       (.I0(\apbi[pwdata] [13]),
        .I1(\r_reg[iforce][3]__0 [12]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [29]),
        .I4(\r[iforce][3][13]_i_2_n_0 ),
        .I5(\r[iforce][3][13]_i_3_n_0 ),
        .O(\r[iforce][3][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][13]_i_2 
       (.I0(\apbi[pirq] [13]),
        .I1(p_0_in8_in),
        .O(\r[iforce][3][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][3][13]_i_3 
       (.I0(\irqi[3][irl] [2]),
        .I1(\irqi[3][irl] [3]),
        .I2(\irqi[3][intack] ),
        .I3(\irqi[3][irl] [0]),
        .I4(\irqi[3][irl] [1]),
        .O(\r[iforce][3][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][14]_i_1 
       (.I0(\apbi[pwdata] [14]),
        .I1(\r_reg[iforce][3]__0 [13]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [30]),
        .I4(\r[iforce][3][14]_i_3_n_0 ),
        .I5(\r[iforce][3][14]_i_4_n_0 ),
        .O(\r[iforce][3][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[iforce][3][14]_i_2 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\r[iforce][3][15]_i_4_n_0 ),
        .O(\r[iforce][3][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][14]_i_3 
       (.I0(\apbi[pirq] [14]),
        .I1(p_0_in6_in),
        .O(\r[iforce][3][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00008000)) 
    \r[iforce][3][14]_i_4 
       (.I0(\irqi[3][irl] [2]),
        .I1(\irqi[3][irl] [3]),
        .I2(\irqi[3][intack] ),
        .I3(\irqi[3][irl] [1]),
        .I4(\irqi[3][irl] [0]),
        .O(\r[iforce][3][14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEA00EAEAEAEAEAEA)) 
    \r[iforce][3][15]_i_1 
       (.I0(\r[iforce][3][15]_i_2_n_0 ),
        .I1(\apbi[pirq] [15]),
        .I2(p_0_in4_in),
        .I3(\r[iforce][3][15]_i_3_n_0 ),
        .I4(\irqi[3][irl] [0]),
        .I5(\irqi[3][irl] [1]),
        .O(\r[iforce][3][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCC0ECCCCCCCCCC)) 
    \r[iforce][3][15]_i_2 
       (.I0(\apbi[pwdata] [15]),
        .I1(\r_reg[iforce][3]__0 [14]),
        .I2(\apbi[pwdata] [31]),
        .I3(\apbi[paddr] [3]),
        .I4(\apbi[paddr] [4]),
        .I5(\r[iforce][3][15]_i_4_n_0 ),
        .O(\r[iforce][3][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7F)) 
    \r[iforce][3][15]_i_3 
       (.I0(\irqi[3][intack] ),
        .I1(\irqi[3][irl] [3]),
        .I2(\irqi[3][irl] [2]),
        .O(\r[iforce][3][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][3][15]_i_4 
       (.I0(\apbi[paddr] [2]),
        .I1(\r[cpurst][0]_i_3_n_0 ),
        .I2(\apbi[paddr] [6]),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [5]),
        .O(\r[iforce][3][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][1]_i_1 
       (.I0(\apbi[pwdata] [1]),
        .I1(\r_reg[iforce][3]__0 [0]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [17]),
        .I4(\r[iforce][3][1]_i_2_n_0 ),
        .I5(\r[iforce][3][1]_i_3_n_0 ),
        .O(\r[iforce][3][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][1]_i_2 
       (.I0(\apbi[pirq] [1]),
        .I1(\r_reg[ibroadcast_n_0_][1] ),
        .O(\r[iforce][3][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][3][1]_i_3 
       (.I0(\irqi[3][irl] [0]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][2]_i_1 
       (.I0(\apbi[pwdata] [2]),
        .I1(\r_reg[iforce][3]__0 [1]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [18]),
        .I4(\r[iforce][3][2]_i_2_n_0 ),
        .I5(\r[iforce][3][2]_i_3_n_0 ),
        .O(\r[iforce][3][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][2]_i_2 
       (.I0(\apbi[pirq] [2]),
        .I1(p_0_in30_in),
        .O(\r[iforce][3][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \r[iforce][3][2]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][3]_i_1 
       (.I0(\apbi[pwdata] [3]),
        .I1(\r_reg[iforce][3]__0 [2]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [19]),
        .I4(\r[iforce][3][3]_i_2_n_0 ),
        .I5(\r[iforce][3][3]_i_3_n_0 ),
        .O(\r[iforce][3][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][3]_i_2 
       (.I0(\apbi[pirq] [3]),
        .I1(p_0_in28_in),
        .O(\r[iforce][3][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000800)) 
    \r[iforce][3][3]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][4]_i_1 
       (.I0(\apbi[pwdata] [4]),
        .I1(\r_reg[iforce][3]__0 [3]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [20]),
        .I4(\r[iforce][3][4]_i_2_n_0 ),
        .I5(\r[iforce][3][4]_i_3_n_0 ),
        .O(\r[iforce][3][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][4]_i_2 
       (.I0(\apbi[pirq] [4]),
        .I1(p_0_in26_in),
        .O(\r[iforce][3][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00100000)) 
    \r[iforce][3][4]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [2]),
        .I3(\irqi[3][irl] [3]),
        .I4(\irqi[3][intack] ),
        .O(\r[iforce][3][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][5]_i_1 
       (.I0(\apbi[pwdata] [5]),
        .I1(\r_reg[iforce][3]__0 [4]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [21]),
        .I4(\r[iforce][3][5]_i_2_n_0 ),
        .I5(\r[iforce][3][5]_i_3_n_0 ),
        .O(\r[iforce][3][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][5]_i_2 
       (.I0(\apbi[pirq] [5]),
        .I1(p_0_in24_in),
        .O(\r[iforce][3][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][3][5]_i_3 
       (.I0(\irqi[3][irl] [0]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [2]),
        .I3(\irqi[3][irl] [3]),
        .I4(\irqi[3][intack] ),
        .O(\r[iforce][3][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][6]_i_1 
       (.I0(\apbi[pwdata] [6]),
        .I1(\r_reg[iforce][3]__0 [5]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [22]),
        .I4(\r[iforce][3][6]_i_2_n_0 ),
        .I5(\r[iforce][3][6]_i_3_n_0 ),
        .O(\r[iforce][3][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][6]_i_2 
       (.I0(\apbi[pirq] [6]),
        .I1(p_0_in22_in),
        .O(\r[iforce][3][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \r[iforce][3][6]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [2]),
        .I3(\irqi[3][irl] [3]),
        .I4(\irqi[3][intack] ),
        .O(\r[iforce][3][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][7]_i_1 
       (.I0(\apbi[pwdata] [7]),
        .I1(\r_reg[iforce][3]__0 [6]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [23]),
        .I4(\r[iforce][3][7]_i_2_n_0 ),
        .I5(\r[iforce][3][7]_i_3_n_0 ),
        .O(\r[iforce][3][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][7]_i_2 
       (.I0(\apbi[pirq] [7]),
        .I1(p_0_in20_in),
        .O(\r[iforce][3][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00800000)) 
    \r[iforce][3][7]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [2]),
        .I3(\irqi[3][irl] [3]),
        .I4(\irqi[3][intack] ),
        .O(\r[iforce][3][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][8]_i_1 
       (.I0(\apbi[pwdata] [8]),
        .I1(\r_reg[iforce][3]__0 [7]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [24]),
        .I4(\r[iforce][3][8]_i_2_n_0 ),
        .I5(\r[iforce][3][8]_i_3_n_0 ),
        .O(\r[iforce][3][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][8]_i_2 
       (.I0(\apbi[pirq] [8]),
        .I1(p_0_in18_in),
        .O(\r[iforce][3][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \r[iforce][3][8]_i_3 
       (.I0(\irqi[3][irl] [1]),
        .I1(\irqi[3][irl] [0]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFFC0CE)) 
    \r[iforce][3][9]_i_1 
       (.I0(\apbi[pwdata] [9]),
        .I1(\r_reg[iforce][3]__0 [8]),
        .I2(\r[iforce][3][14]_i_2_n_0 ),
        .I3(\apbi[pwdata] [25]),
        .I4(\r[iforce][3][9]_i_2_n_0 ),
        .I5(\r[iforce][3][9]_i_3_n_0 ),
        .O(\r[iforce][3][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \r[iforce][3][9]_i_2 
       (.I0(\apbi[pirq] [9]),
        .I1(p_0_in16_in),
        .O(\r[iforce][3][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \r[iforce][3][9]_i_3 
       (.I0(\irqi[3][irl] [0]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [3]),
        .I3(\irqi[3][intack] ),
        .I4(\irqi[3][irl] [2]),
        .O(\r[iforce][3][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[ilevel][15]_i_1 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\r[cpurst][0]_i_3_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [2]),
        .I5(\apbi[paddr] [6]),
        .O(\v[ilevel] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \r[imask][0][15]_i_1 
       (.I0(\apbi[paddr] [4]),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [6]),
        .I3(\apbi[paddr] [5]),
        .I4(\r[imask][0][15]_i_2_n_0 ),
        .O(\v[imask][0] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    \r[imask][0][15]_i_2 
       (.I0(\apbi[pwrite] ),
        .I1(apbi[2]),
        .I2(\apbi[penable] ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [2]),
        .O(\r[imask][0][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00400000)) 
    \r[imask][1][15]_i_1 
       (.I0(\r[cpurst][0]_i_3_n_0 ),
        .I1(\apbi[paddr] [2]),
        .I2(\r[imask][1][15]_i_2_n_0 ),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [6]),
        .O(\v[imask][1] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \r[imask][1][15]_i_2 
       (.I0(\apbi[paddr] [3]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [5]),
        .O(\r[imask][1][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    \r[imask][2][15]_i_1 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [7]),
        .I2(\r[cpurst][0]_i_3_n_0 ),
        .I3(\apbi[paddr] [6]),
        .I4(\r[imask][2][15]_i_2_n_0 ),
        .O(\v[imask][2] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \r[imask][2][15]_i_2 
       (.I0(\apbi[paddr] [5]),
        .I1(\apbi[paddr] [3]),
        .I2(\apbi[paddr] [4]),
        .O(\r[imask][2][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \r[imask][3][15]_i_1 
       (.I0(\r[forceerr][0]_i_3_n_0 ),
        .I1(\apbi[paddr] [6]),
        .I2(\apbi[paddr] [5]),
        .I3(\apbi[paddr] [7]),
        .I4(\apbi[paddr] [4]),
        .I5(\apbi[paddr] [2]),
        .O(\v[imask][3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022202220220000)) 
    \r[ipend][10]_i_1 
       (.I0(\r[ipend][10]_i_2_n_0 ),
        .I1(\r[ipend][10]_i_3_n_0 ),
        .I2(\r_reg[iforce][1]__0 [9]),
        .I3(\r[iforce][1][10]_i_2_n_0 ),
        .I4(\r[ipend][10]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [9]),
        .O(\r[ipend][10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][10]_i_2 
       (.I0(p_0_in14_in),
        .I1(\apbi[pirq] [10]),
        .I2(\apbi[pwdata] [10]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[10]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[ipend][10]_i_3 
       (.I0(\r_reg[iforce][3]__0 [9]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [0]),
        .I3(\r[ipend][10]_i_5_n_0 ),
        .I4(\r_reg[iforce][2]__0 [9]),
        .I5(\r[iforce][2][10]_i_2_n_0 ),
        .O(\r[ipend][10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFDFFF)) 
    \r[ipend][10]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r[ipend][10]_i_5 
       (.I0(\irqi[3][irl] [2]),
        .I1(\irqi[3][intack] ),
        .I2(\irqi[3][irl] [3]),
        .O(\r[ipend][10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022202220220000)) 
    \r[ipend][11]_i_1 
       (.I0(\r[ipend][11]_i_2_n_0 ),
        .I1(\r[ipend][11]_i_3_n_0 ),
        .I2(\r_reg[iforce][1]__0 [10]),
        .I3(\r[iforce][1][11]_i_2_n_0 ),
        .I4(\r[ipend][11]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [10]),
        .O(\r[ipend][11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][11]_i_2 
       (.I0(p_0_in12_in),
        .I1(\apbi[pirq] [11]),
        .I2(\apbi[pwdata] [11]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[11]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \r[ipend][11]_i_3 
       (.I0(\r_reg[iforce][2]__0 [10]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [0]),
        .I3(\r[ipend][11]_i_5_n_0 ),
        .I4(\r_reg[iforce][3]__0 [10]),
        .I5(\r[iforce][3][11]_i_3_n_0 ),
        .O(\r[ipend][11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \r[ipend][11]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \r[ipend][11]_i_5 
       (.I0(\irqi[2][irl] [2]),
        .I1(\irqi[2][intack] ),
        .I2(\irqi[2][irl] [3]),
        .O(\r[ipend][11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220000022202220)) 
    \r[ipend][12]_i_1 
       (.I0(\r[ipend][12]_i_2_n_0 ),
        .I1(\r[ipend][12]_i_3_n_0 ),
        .I2(\r[ipend][12]_i_4_n_0 ),
        .I3(\r_reg[iforce][0]__0 [11]),
        .I4(\r_reg[iforce][1]__0 [11]),
        .I5(\r[iforce][1][12]_i_2_n_0 ),
        .O(\r[ipend][12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][12]_i_2 
       (.I0(p_0_in10_in),
        .I1(\apbi[pirq] [12]),
        .I2(\apbi[pwdata] [12]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[12]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001FFFF00010001)) 
    \r[ipend][12]_i_3 
       (.I0(\r_reg[iforce][2]__0 [11]),
        .I1(\r[iforce][2][15]_i_3_n_0 ),
        .I2(\irqi[2][irl] [1]),
        .I3(\irqi[2][irl] [0]),
        .I4(\r_reg[iforce][3]__0 [11]),
        .I5(\r[iforce][3][12]_i_3_n_0 ),
        .O(\r[ipend][12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFF7F)) 
    \r[ipend][12]_i_4 
       (.I0(\irqi[0][irl] [2]),
        .I1(\irqi[0][irl] [3]),
        .I2(irqi),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .O(\r[ipend][12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220000022202220)) 
    \r[ipend][13]_i_1 
       (.I0(\r[ipend][13]_i_2_n_0 ),
        .I1(\r[ipend][13]_i_3_n_0 ),
        .I2(\r[ipend][13]_i_4_n_0 ),
        .I3(\r_reg[iforce][0]__0 [12]),
        .I4(\r_reg[iforce][1]__0 [12]),
        .I5(\r[iforce][1][13]_i_2_n_0 ),
        .O(\r[ipend][13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][13]_i_2 
       (.I0(p_0_in8_in),
        .I1(\apbi[pirq] [13]),
        .I2(\apbi[pwdata] [13]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[13]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100010)) 
    \r[ipend][13]_i_3 
       (.I0(\r_reg[iforce][2]__0 [12]),
        .I1(\r[iforce][2][15]_i_3_n_0 ),
        .I2(\irqi[2][irl] [0]),
        .I3(\irqi[2][irl] [1]),
        .I4(\r_reg[iforce][3]__0 [12]),
        .I5(\r[iforce][3][13]_i_3_n_0 ),
        .O(\r[ipend][13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \r[ipend][13]_i_4 
       (.I0(\irqi[0][irl] [2]),
        .I1(\irqi[0][irl] [3]),
        .I2(irqi),
        .I3(\irqi[0][irl] [0]),
        .I4(\irqi[0][irl] [1]),
        .O(\r[ipend][13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022202220220000)) 
    \r[ipend][14]_i_1 
       (.I0(\r[ipend][14]_i_2_n_0 ),
        .I1(\r[ipend][14]_i_3_n_0 ),
        .I2(\r_reg[iforce][1]__0 [13]),
        .I3(\r[iforce][1][14]_i_2_n_0 ),
        .I4(\r[ipend][14]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [13]),
        .O(\r[ipend][14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][14]_i_2 
       (.I0(p_0_in6_in),
        .I1(\apbi[pirq] [14]),
        .I2(\apbi[pwdata] [14]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[14]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100010)) 
    \r[ipend][14]_i_3 
       (.I0(\r_reg[iforce][2]__0 [13]),
        .I1(\r[iforce][2][15]_i_3_n_0 ),
        .I2(\irqi[2][irl] [1]),
        .I3(\irqi[2][irl] [0]),
        .I4(\r_reg[iforce][3]__0 [13]),
        .I5(\r[iforce][3][14]_i_4_n_0 ),
        .O(\r[ipend][14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF7FFF)) 
    \r[ipend][14]_i_4 
       (.I0(\irqi[0][irl] [2]),
        .I1(\irqi[0][irl] [3]),
        .I2(irqi),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .O(\r[ipend][14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    \r[ipend][15]_i_1 
       (.I0(\r[ipend][15]_i_2_n_0 ),
        .I1(\r[ipend][15]_i_3_n_0 ),
        .I2(\r_reg[iforce][2]__0 [14]),
        .I3(\r[ipend][15]_i_4_n_0 ),
        .I4(\r_reg[iforce][1]__0 [14]),
        .I5(\r[iforce][1][15]_i_4_n_0 ),
        .O(\r[ipend][15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][15]_i_2 
       (.I0(p_0_in4_in),
        .I1(\apbi[pirq] [15]),
        .I2(\apbi[pwdata] [15]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[15]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h004000400040FFFF)) 
    \r[ipend][15]_i_3 
       (.I0(\r_reg[iforce][3]__0 [14]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [0]),
        .I3(\r[iforce][3][15]_i_3_n_0 ),
        .I4(\r[ipend][15]_i_6_n_0 ),
        .I5(\r_reg[iforce][0]__0 [14]),
        .O(\r[ipend][15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \r[ipend][15]_i_4 
       (.I0(\irqi[2][irl] [1]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [2]),
        .I3(\irqi[2][irl] [3]),
        .I4(\irqi[2][intack] ),
        .O(\r[ipend][15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFD)) 
    \r[ipend][15]_i_5 
       (.I0(\apbi[paddr] [2]),
        .I1(\apbi[paddr] [4]),
        .I2(\apbi[paddr] [7]),
        .I3(\r[cpurst][0]_i_3_n_0 ),
        .I4(\apbi[paddr] [6]),
        .O(\r[ipend][15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h7FFFFFFF)) 
    \r[ipend][15]_i_6 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [3]),
        .I4(irqi),
        .O(\r[ipend][15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220000022202220)) 
    \r[ipend][1]_i_1 
       (.I0(\r[ipend][1]_i_2_n_0 ),
        .I1(\r[ipend][1]_i_3_n_0 ),
        .I2(\r[ipend][1]_i_4_n_0 ),
        .I3(\r_reg[iforce][0]__0 [0]),
        .I4(\r_reg[iforce][1]__0 [0]),
        .I5(\r[iforce][1][1]_i_2_n_0 ),
        .O(\r[ipend][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][1]_i_2 
       (.I0(\r_reg[ibroadcast_n_0_][1] ),
        .I1(\apbi[pirq] [1]),
        .I2(\apbi[pwdata] [1]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[1]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[ipend][1]_i_3 
       (.I0(\r_reg[iforce][2]__0 [0]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [1]),
        .I3(\r[ipend][3]_i_5_n_0 ),
        .I4(\r_reg[iforce][3]__0 [0]),
        .I5(\r[iforce][3][1]_i_3_n_0 ),
        .O(\r[ipend][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFDFF)) 
    \r[ipend][1]_i_4 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022202220220000)) 
    \r[ipend][2]_i_1 
       (.I0(\r[ipend][2]_i_2_n_0 ),
        .I1(\r[ipend][2]_i_3_n_0 ),
        .I2(\r_reg[iforce][1]__0 [1]),
        .I3(\r[iforce][1][2]_i_2_n_0 ),
        .I4(\r[ipend][2]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [1]),
        .O(\r[ipend][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][2]_i_2 
       (.I0(p_0_in30_in),
        .I1(\apbi[pirq] [2]),
        .I2(\apbi[pwdata] [2]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[2]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[ipend][2]_i_3 
       (.I0(\r_reg[iforce][2]__0 [1]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [0]),
        .I3(\r[ipend][3]_i_5_n_0 ),
        .I4(\r_reg[iforce][3]__0 [1]),
        .I5(\r[iforce][3][2]_i_3_n_0 ),
        .O(\r[ipend][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFDFF)) 
    \r[ipend][2]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022202220220000)) 
    \r[ipend][3]_i_1 
       (.I0(\r[ipend][3]_i_2_n_0 ),
        .I1(\r[ipend][3]_i_3_n_0 ),
        .I2(\r_reg[iforce][1]__0 [2]),
        .I3(\r[iforce][1][3]_i_2_n_0 ),
        .I4(\r[ipend][3]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [2]),
        .O(\r[ipend][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][3]_i_2 
       (.I0(p_0_in28_in),
        .I1(\apbi[pirq] [3]),
        .I2(\apbi[pwdata] [3]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[3]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \r[ipend][3]_i_3 
       (.I0(\r_reg[iforce][2]__0 [2]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [0]),
        .I3(\r[ipend][3]_i_5_n_0 ),
        .I4(\r_reg[iforce][3]__0 [2]),
        .I5(\r[iforce][3][3]_i_3_n_0 ),
        .O(\r[ipend][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF7FF)) 
    \r[ipend][3]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \r[ipend][3]_i_5 
       (.I0(\irqi[2][irl] [2]),
        .I1(\irqi[2][intack] ),
        .I2(\irqi[2][irl] [3]),
        .O(\r[ipend][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    \r[ipend][4]_i_1 
       (.I0(\r[ipend][4]_i_2_n_0 ),
        .I1(\r[ipend][4]_i_3_n_0 ),
        .I2(\r_reg[iforce][2]__0 [3]),
        .I3(\r[iforce][2][4]_i_2_n_0 ),
        .I4(\r_reg[iforce][1]__0 [3]),
        .I5(\r[iforce][1][4]_i_2_n_0 ),
        .O(\r[ipend][4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][4]_i_2 
       (.I0(p_0_in26_in),
        .I1(\apbi[pirq] [4]),
        .I2(\apbi[pwdata] [4]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[4]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000100010001FFFF)) 
    \r[ipend][4]_i_3 
       (.I0(\r_reg[iforce][3]__0 [3]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [0]),
        .I3(\r[ipend][7]_i_5_n_0 ),
        .I4(\r[ipend][4]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [3]),
        .O(\r[ipend][4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFDF)) 
    \r[ipend][4]_i_4 
       (.I0(\irqi[0][irl] [2]),
        .I1(\irqi[0][irl] [3]),
        .I2(irqi),
        .I3(\irqi[0][irl] [1]),
        .I4(\irqi[0][irl] [0]),
        .O(\r[ipend][4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    \r[ipend][5]_i_1 
       (.I0(\r[ipend][5]_i_2_n_0 ),
        .I1(\r[ipend][5]_i_3_n_0 ),
        .I2(\r_reg[iforce][3]__0 [4]),
        .I3(\r[iforce][3][5]_i_3_n_0 ),
        .I4(\r_reg[iforce][1]__0 [4]),
        .I5(\r[iforce][1][5]_i_2_n_0 ),
        .O(\r[ipend][5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][5]_i_2 
       (.I0(p_0_in24_in),
        .I1(\apbi[pirq] [5]),
        .I2(\apbi[pwdata] [5]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[5]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000400040004FFFF)) 
    \r[ipend][5]_i_3 
       (.I0(\r_reg[iforce][2]__0 [4]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [1]),
        .I3(\r[ipend][6]_i_5_n_0 ),
        .I4(\r[ipend][5]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [4]),
        .O(\r[ipend][5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \r[ipend][5]_i_4 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [3]),
        .I4(irqi),
        .O(\r[ipend][5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220000022202220)) 
    \r[ipend][6]_i_1 
       (.I0(\r[ipend][6]_i_2_n_0 ),
        .I1(\r[ipend][6]_i_3_n_0 ),
        .I2(\r[ipend][6]_i_4_n_0 ),
        .I3(\r_reg[iforce][0]__0 [5]),
        .I4(\r_reg[iforce][1]__0 [5]),
        .I5(\r[iforce][1][6]_i_2_n_0 ),
        .O(\r[ipend][6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][6]_i_2 
       (.I0(p_0_in22_in),
        .I1(\apbi[pirq] [6]),
        .I2(\apbi[pwdata] [6]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[6]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040004)) 
    \r[ipend][6]_i_3 
       (.I0(\r_reg[iforce][2]__0 [5]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [0]),
        .I3(\r[ipend][6]_i_5_n_0 ),
        .I4(\r_reg[iforce][3]__0 [5]),
        .I5(\r[iforce][3][6]_i_3_n_0 ),
        .O(\r[ipend][6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFDFFFFF)) 
    \r[ipend][6]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [3]),
        .I4(irqi),
        .O(\r[ipend][6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[ipend][6]_i_5 
       (.I0(\irqi[2][intack] ),
        .I1(\irqi[2][irl] [3]),
        .I2(\irqi[2][irl] [2]),
        .O(\r[ipend][6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2220000022202220)) 
    \r[ipend][7]_i_1 
       (.I0(\r[ipend][7]_i_2_n_0 ),
        .I1(\r[ipend][7]_i_3_n_0 ),
        .I2(\r[ipend][7]_i_4_n_0 ),
        .I3(\r_reg[iforce][0]__0 [6]),
        .I4(\r_reg[iforce][1]__0 [6]),
        .I5(\r[iforce][1][7]_i_2_n_0 ),
        .O(\r[ipend][7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][7]_i_2 
       (.I0(p_0_in20_in),
        .I1(\apbi[pirq] [7]),
        .I2(\apbi[pwdata] [7]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[7]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0040FFFF00400040)) 
    \r[ipend][7]_i_3 
       (.I0(\r_reg[iforce][3]__0 [6]),
        .I1(\irqi[3][irl] [1]),
        .I2(\irqi[3][irl] [0]),
        .I3(\r[ipend][7]_i_5_n_0 ),
        .I4(\r_reg[iforce][2]__0 [6]),
        .I5(\r[iforce][2][7]_i_2_n_0 ),
        .O(\r[ipend][7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF7FFFFF)) 
    \r[ipend][7]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [2]),
        .I3(\irqi[0][irl] [3]),
        .I4(irqi),
        .O(\r[ipend][7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hDF)) 
    \r[ipend][7]_i_5 
       (.I0(\irqi[3][intack] ),
        .I1(\irqi[3][irl] [3]),
        .I2(\irqi[3][irl] [2]),
        .O(\r[ipend][7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    \r[ipend][8]_i_1 
       (.I0(\r[ipend][8]_i_2_n_0 ),
        .I1(\r[ipend][8]_i_3_n_0 ),
        .I2(\r_reg[iforce][3]__0 [7]),
        .I3(\r[iforce][3][8]_i_3_n_0 ),
        .I4(\r_reg[iforce][1]__0 [7]),
        .I5(\r[iforce][1][8]_i_2_n_0 ),
        .O(\r[ipend][8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][8]_i_2 
       (.I0(p_0_in18_in),
        .I1(\apbi[pirq] [8]),
        .I2(\apbi[pwdata] [8]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[8]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001FFFF00010001)) 
    \r[ipend][8]_i_3 
       (.I0(\r_reg[iforce][2]__0 [7]),
        .I1(\irqi[2][irl] [1]),
        .I2(\irqi[2][irl] [0]),
        .I3(\r[ipend][11]_i_5_n_0 ),
        .I4(\r_reg[iforce][0]__0 [7]),
        .I5(\r[ipend][8]_i_4_n_0 ),
        .O(\r[ipend][8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \r[ipend][8]_i_4 
       (.I0(\irqi[0][irl] [1]),
        .I1(\irqi[0][irl] [0]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2022000020222022)) 
    \r[ipend][9]_i_1 
       (.I0(\r[ipend][9]_i_2_n_0 ),
        .I1(\r[ipend][9]_i_3_n_0 ),
        .I2(\r_reg[iforce][3]__0 [8]),
        .I3(\r[iforce][3][9]_i_3_n_0 ),
        .I4(\r_reg[iforce][1]__0 [8]),
        .I5(\r[iforce][1][9]_i_2_n_0 ),
        .O(\r[ipend][9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF44444FF444F4)) 
    \r[ipend][9]_i_2 
       (.I0(p_0_in16_in),
        .I1(\apbi[pirq] [9]),
        .I2(\apbi[pwdata] [9]),
        .I3(\apbi[paddr] [3]),
        .I4(p_5_in[9]),
        .I5(\r[ipend][15]_i_5_n_0 ),
        .O(\r[ipend][9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000400040004FFFF)) 
    \r[ipend][9]_i_3 
       (.I0(\r_reg[iforce][2]__0 [8]),
        .I1(\irqi[2][irl] [0]),
        .I2(\irqi[2][irl] [1]),
        .I3(\r[ipend][11]_i_5_n_0 ),
        .I4(\r[ipend][9]_i_4_n_0 ),
        .I5(\r_reg[iforce][0]__0 [8]),
        .O(\r[ipend][9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFDFFF)) 
    \r[ipend][9]_i_4 
       (.I0(\irqi[0][irl] [0]),
        .I1(\irqi[0][irl] [1]),
        .I2(\irqi[0][irl] [3]),
        .I3(irqi),
        .I4(\irqi[0][irl] [2]),
        .O(\r[ipend][9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFAFAFACA0A0A0AC)) 
    \r[irl][0][0]_i_1 
       (.I0(\r[irl][0][0]_i_2_n_0 ),
        .I1(\r[irl][0][0]_i_3_n_0 ),
        .I2(\r[irl][0][2]_i_6_n_0 ),
        .I3(\r[irl][0][0]_i_4_n_0 ),
        .I4(\r[irl][0][3]_i_4_n_0 ),
        .I5(\r[irl][0][0]_i_5_n_0 ),
        .O(\r[irl][0][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF000C00FF000E00)) 
    \r[irl][0][0]_i_10 
       (.I0(\r[irl][0][3]_i_15_n_0 ),
        .I1(\r[irl][0][2]_i_10_n_0 ),
        .I2(\r[irl][0][2]_i_9_n_0 ),
        .I3(\r[irl][0][2]_i_8_n_0 ),
        .I4(\r[irl][0][2]_i_7_n_0 ),
        .I5(\r[irl][0][3]_i_16_n_0 ),
        .O(\r[irl][0][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFF4544)) 
    \r[irl][0][0]_i_11 
       (.I0(\r[irl][0][3]_i_13_n_0 ),
        .I1(\r[irl][0][2]_i_21_n_0 ),
        .I2(\r[irl][0][2]_i_17_n_0 ),
        .I3(\r[irl][0][0]_i_12_n_0 ),
        .I4(\r[irl][0][1]_i_11_n_0 ),
        .I5(\r[irl][0][3]_i_21_n_0 ),
        .O(\r[irl][0][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][0]_i_12 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][0]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][0]__0 [4]),
        .O(\r[irl][0][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF004F00FF)) 
    \r[irl][0][0]_i_2 
       (.I0(\r[irl][0][2]_i_19_n_0 ),
        .I1(p_6_in[3]),
        .I2(\r[irl][0][3]_i_11_n_0 ),
        .I3(\r[irl][0][0]_i_6_n_0 ),
        .I4(\r[irl][0][3]_i_10_n_0 ),
        .I5(\r[irl][0][3]_i_9_n_0 ),
        .O(\r[irl][0][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][0]_i_3 
       (.I0(p_6_in[1]),
        .I1(\r_reg[iforce][0]__0 [0]),
        .I2(p_5_in[1]),
        .I3(\r_reg[imask][0]__0 [0]),
        .O(\r[irl][0][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEFEFEFF)) 
    \r[irl][0][0]_i_4 
       (.I0(\r[irl][0][0]_i_7_n_0 ),
        .I1(\r[irl][0][2]_i_18_n_0 ),
        .I2(\r[irl][0][2]_i_17_n_0 ),
        .I3(\r[irl][0][0]_i_8_n_0 ),
        .I4(p_6_in[2]),
        .O(\r[irl][0][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCCCCCCCCCCCCC8A)) 
    \r[irl][0][0]_i_5 
       (.I0(\r[irl][0][0]_i_7_n_0 ),
        .I1(\r[irl][0][0]_i_9_n_0 ),
        .I2(\r[irl][0][2]_i_16_n_0 ),
        .I3(\r[irl][0][2]_i_17_n_0 ),
        .I4(\r[irl][0][2]_i_18_n_0 ),
        .I5(\r[irl][0][3]_i_4_n_0 ),
        .O(\r[irl][0][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0FFF0F0F0F2)) 
    \r[irl][0][0]_i_6 
       (.I0(\r[irl][0][1]_i_6_n_0 ),
        .I1(\r[irl][0][3]_i_18_n_0 ),
        .I2(\r[irl][0][0]_i_10_n_0 ),
        .I3(\r[irl][0][3]_i_17_n_0 ),
        .I4(\r[irl][0][3]_i_6_n_0 ),
        .I5(\r[irl][0][3]_i_5_n_0 ),
        .O(\r[irl][0][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00A8)) 
    \r[irl][0][0]_i_7 
       (.I0(\r_reg[imask][0]__0 [2]),
        .I1(p_5_in[3]),
        .I2(\r_reg[iforce][0]__0 [2]),
        .I3(p_6_in[3]),
        .I4(\r[irl][0][2]_i_16_n_0 ),
        .O(\r[irl][0][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][0][0]_i_8 
       (.I0(\r_reg[imask][0]__0 [1]),
        .I1(p_5_in[2]),
        .I2(\r_reg[iforce][0]__0 [1]),
        .O(\r[irl][0][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFF0F0F0FFF0FE)) 
    \r[irl][0][0]_i_9 
       (.I0(\r[irl][0][0]_i_11_n_0 ),
        .I1(\r[irl][0][3]_i_22_n_0 ),
        .I2(\r[irl][0][2]_i_12_n_0 ),
        .I3(\r[irl][0][2]_i_13_n_0 ),
        .I4(\r[irl][0][2]_i_14_n_0 ),
        .I5(\r[irl][0][2]_i_15_n_0 ),
        .O(\r[irl][0][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hD0FFD0D0D0FFD0FF)) 
    \r[irl][0][1]_i_1 
       (.I0(\r[irl][0][2]_i_3_n_0 ),
        .I1(\r[irl][0][1]_i_2_n_0 ),
        .I2(\r[irl][0][1]_i_3_n_0 ),
        .I3(\r[irl][0][3]_i_3_n_0 ),
        .I4(\r[irl][0][1]_i_4_n_0 ),
        .I5(\r[irl][0][2]_i_5_n_0 ),
        .O(\r[irl][0][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][0][1]_i_10 
       (.I0(\r_reg[imask][0]__0 [13]),
        .I1(p_5_in[14]),
        .I2(\r_reg[iforce][0]__0 [13]),
        .I3(p_6_in[14]),
        .I4(\r[irl][0][2]_i_12_n_0 ),
        .O(\r[irl][0][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][1]_i_11 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][0]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][0]__0 [8]),
        .O(\r[irl][0][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][0][1]_i_12 
       (.I0(\r_reg[imask][0]__0 [10]),
        .I1(p_5_in[11]),
        .I2(\r_reg[iforce][0]__0 [10]),
        .O(\r[irl][0][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA800)) 
    \r[irl][0][1]_i_13 
       (.I0(\r_reg[imask][0]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][0]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][0][2]_i_9_n_0 ),
        .O(\r[irl][0][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000777F)) 
    \r[irl][0][1]_i_14 
       (.I0(p_6_in[15]),
        .I1(\r_reg[imask][0]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[iforce][0]__0 [14]),
        .I4(\r[irl][0][2]_i_7_n_0 ),
        .O(\r[irl][0][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00F4F4)) 
    \r[irl][0][1]_i_2 
       (.I0(\r[irl][0][1]_i_5_n_0 ),
        .I1(p_6_in[7]),
        .I2(\r[irl][0][1]_i_6_n_0 ),
        .I3(\r[irl][0][1]_i_7_n_0 ),
        .I4(\r[irl][0][3]_i_2_n_0 ),
        .O(\r[irl][0][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF2FF)) 
    \r[irl][0][1]_i_3 
       (.I0(p_6_in[3]),
        .I1(\r[irl][0][2]_i_19_n_0 ),
        .I2(\r[irl][0][3]_i_9_n_0 ),
        .I3(\r[irl][0][3]_i_10_n_0 ),
        .I4(\r[irl][0][3]_i_11_n_0 ),
        .O(\r[irl][0][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC0CCC0CCC0CCD1DD)) 
    \r[irl][0][1]_i_4 
       (.I0(\r[irl][0][1]_i_8_n_0 ),
        .I1(\r[irl][0][3]_i_14_n_0 ),
        .I2(\r[irl][0][1]_i_9_n_0 ),
        .I3(\r[irl][0][1]_i_10_n_0 ),
        .I4(\r[irl][0][3]_i_13_n_0 ),
        .I5(\r[irl][0][1]_i_11_n_0 ),
        .O(\r[irl][0][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][0][1]_i_5 
       (.I0(\r_reg[imask][0]__0 [6]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][0]__0 [6]),
        .O(\r[irl][0][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][1]_i_6 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][0]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][0]__0 [5]),
        .O(\r[irl][0][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00F4FFFF)) 
    \r[irl][0][1]_i_7 
       (.I0(\r[irl][0][1]_i_12_n_0 ),
        .I1(p_6_in[11]),
        .I2(\r[irl][0][3]_i_15_n_0 ),
        .I3(\r[irl][0][1]_i_13_n_0 ),
        .I4(\r[irl][0][1]_i_14_n_0 ),
        .O(\r[irl][0][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551115)) 
    \r[irl][0][1]_i_8 
       (.I0(\r[irl][0][2]_i_17_n_0 ),
        .I1(\r_reg[imask][0]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[iforce][0]__0 [6]),
        .I4(p_6_in[7]),
        .O(\r[irl][0][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][0][1]_i_9 
       (.I0(\r_reg[imask][0]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][0]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][0][2]_i_14_n_0 ),
        .O(\r[irl][0][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7070707070FF7070)) 
    \r[irl][0][2]_i_1 
       (.I0(\r[irl][0][2]_i_2_n_0 ),
        .I1(\r[irl][0][3]_i_2_n_0 ),
        .I2(\r[irl][0][2]_i_3_n_0 ),
        .I3(\r[irl][0][2]_i_4_n_0 ),
        .I4(\r[irl][0][2]_i_5_n_0 ),
        .I5(\r[irl][0][2]_i_6_n_0 ),
        .O(\r[irl][0][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][2]_i_10 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][0]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][0]__0 [11]),
        .O(\r[irl][0][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    \r[irl][0][2]_i_11 
       (.I0(\r[irl][0][1]_i_6_n_0 ),
        .I1(\r[irl][0][3]_i_18_n_0 ),
        .I2(\r[irl][0][3]_i_5_n_0 ),
        .I3(p_6_in[9]),
        .I4(\r[irl][0][2]_i_20_n_0 ),
        .I5(\r[irl][0][3]_i_6_n_0 ),
        .O(\r[irl][0][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_12 
       (.I0(p_6_in[15]),
        .I1(\r_reg[iforce][0]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[imask][0]__0 [14]),
        .O(\r[irl][0][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_13 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][0]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][0]__0 [13]),
        .O(\r[irl][0][2]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_14 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][0]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][0]__0 [12]),
        .O(\r[irl][0][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_15 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][0]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][0]__0 [11]),
        .O(\r[irl][0][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_16 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][0]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][0]__0 [3]),
        .O(\r[irl][0][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_17 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][0]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][0]__0 [5]),
        .O(\r[irl][0][2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAEEEA)) 
    \r[irl][0][2]_i_18 
       (.I0(\r[irl][0][2]_i_21_n_0 ),
        .I1(\r_reg[imask][0]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[iforce][0]__0 [4]),
        .I4(p_6_in[5]),
        .O(\r[irl][0][2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][0][2]_i_19 
       (.I0(\r_reg[imask][0]__0 [2]),
        .I1(p_5_in[3]),
        .I2(\r_reg[iforce][0]__0 [2]),
        .O(\r[irl][0][2]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \r[irl][0][2]_i_2 
       (.I0(\r[irl][0][2]_i_7_n_0 ),
        .I1(\r[irl][0][2]_i_8_n_0 ),
        .I2(\r[irl][0][2]_i_9_n_0 ),
        .I3(\r[irl][0][2]_i_10_n_0 ),
        .O(\r[irl][0][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][0][2]_i_20 
       (.I0(\r_reg[imask][0]__0 [8]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][0]__0 [8]),
        .O(\r[irl][0][2]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][2]_i_21 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][0]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][0]__0 [6]),
        .O(\r[irl][0][2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][0][2]_i_3 
       (.I0(\r[irl][0][3]_i_9_n_0 ),
        .I1(p_6_in[5]),
        .I2(\r_reg[iforce][0]__0 [4]),
        .I3(p_5_in[5]),
        .I4(\r_reg[imask][0]__0 [4]),
        .I5(\r[irl][0][2]_i_11_n_0 ),
        .O(\r[irl][0][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \r[irl][0][2]_i_4 
       (.I0(\r[irl][0][2]_i_12_n_0 ),
        .I1(\r[irl][0][2]_i_13_n_0 ),
        .I2(\r[irl][0][2]_i_14_n_0 ),
        .I3(\r[irl][0][2]_i_15_n_0 ),
        .I4(\r[irl][0][3]_i_4_n_0 ),
        .O(\r[irl][0][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \r[irl][0][2]_i_5 
       (.I0(\r[irl][0][2]_i_16_n_0 ),
        .I1(\r[irl][0][2]_i_17_n_0 ),
        .I2(\r[irl][0][2]_i_18_n_0 ),
        .I3(\r[irl][0][3]_i_4_n_0 ),
        .O(\r[irl][0][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFBFFFBFB)) 
    \r[irl][0][2]_i_6 
       (.I0(\r[irl][0][3]_i_11_n_0 ),
        .I1(\r[irl][0][3]_i_10_n_0 ),
        .I2(\r[irl][0][3]_i_9_n_0 ),
        .I3(\r[irl][0][2]_i_19_n_0 ),
        .I4(p_6_in[3]),
        .I5(\r[irl][0][3]_i_7_n_0 ),
        .O(\r[irl][0][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][2]_i_7 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][0]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][0]__0 [13]),
        .O(\r[irl][0][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1FFF)) 
    \r[irl][0][2]_i_8 
       (.I0(\r_reg[iforce][0]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[imask][0]__0 [14]),
        .I3(p_6_in[15]),
        .O(\r[irl][0][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][2]_i_9 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][0]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][0]__0 [12]),
        .O(\r[irl][0][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \r[irl][0][3]_i_1 
       (.I0(\r[irl][0][3]_i_2_n_0 ),
        .I1(\r[irl][0][3]_i_3_n_0 ),
        .I2(\r[irl][0][3]_i_4_n_0 ),
        .O(\r[irl][0][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[irl][0][3]_i_10 
       (.I0(\r[irl][0][3]_i_6_n_0 ),
        .I1(\r[irl][0][3]_i_17_n_0 ),
        .I2(\r[irl][0][3]_i_5_n_0 ),
        .I3(\r[irl][0][3]_i_18_n_0 ),
        .I4(\r[irl][0][1]_i_6_n_0 ),
        .I5(\r[irl][0][3]_i_19_n_0 ),
        .O(\r[irl][0][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_11 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][0]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][0]__0 [1]),
        .O(\r[irl][0][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[irl][0][3]_i_12 
       (.I0(\r[irl][0][1]_i_11_n_0 ),
        .I1(\r[irl][0][3]_i_14_n_0 ),
        .I2(\r[irl][0][3]_i_13_n_0 ),
        .I3(\r[irl][0][3]_i_20_n_0 ),
        .I4(\r[irl][0][2]_i_18_n_0 ),
        .I5(\r[irl][0][0]_i_7_n_0 ),
        .O(\r[irl][0][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][3]_i_13 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][0]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][0]__0 [7]),
        .O(\r[irl][0][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \r[irl][0][3]_i_14 
       (.I0(\r[irl][0][3]_i_21_n_0 ),
        .I1(\r[irl][0][3]_i_22_n_0 ),
        .I2(\r[irl][0][2]_i_12_n_0 ),
        .I3(\r[irl][0][2]_i_13_n_0 ),
        .I4(\r[irl][0][2]_i_14_n_0 ),
        .I5(\r[irl][0][2]_i_15_n_0 ),
        .O(\r[irl][0][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_15 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][0]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][0]__0 [9]),
        .O(\r[irl][0][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_16 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][0]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][0]__0 [10]),
        .O(\r[irl][0][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_17 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][0]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][0]__0 [8]),
        .O(\r[irl][0][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_18 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][0]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][0]__0 [6]),
        .O(\r[irl][0][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_19 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][0]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][0]__0 [4]),
        .O(\r[irl][0][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][0][3]_i_2 
       (.I0(\r[irl][0][3]_i_5_n_0 ),
        .I1(p_6_in[9]),
        .I2(\r_reg[iforce][0]__0 [8]),
        .I3(p_5_in[9]),
        .I4(\r_reg[imask][0]__0 [8]),
        .I5(\r[irl][0][3]_i_6_n_0 ),
        .O(\r[irl][0][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAEEEA)) 
    \r[irl][0][3]_i_20 
       (.I0(\r[irl][0][2]_i_17_n_0 ),
        .I1(\r_reg[imask][0]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[iforce][0]__0 [1]),
        .I4(p_6_in[2]),
        .O(\r[irl][0][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][3]_i_21 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][0]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][0]__0 [9]),
        .O(\r[irl][0][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][0][3]_i_22 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][0]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][0]__0 [10]),
        .O(\r[irl][0][3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \r[irl][0][3]_i_3 
       (.I0(\r[irl][0][3]_i_7_n_0 ),
        .I1(\r[irl][0][3]_i_8_n_0 ),
        .I2(\r[irl][0][3]_i_9_n_0 ),
        .I3(\r[irl][0][3]_i_10_n_0 ),
        .I4(\r[irl][0][3]_i_11_n_0 ),
        .I5(\r[irl][0][3]_i_12_n_0 ),
        .O(\r[irl][0][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEFEFEEEEEEEEEE)) 
    \r[irl][0][3]_i_4 
       (.I0(\r[irl][0][3]_i_13_n_0 ),
        .I1(\r[irl][0][3]_i_14_n_0 ),
        .I2(p_6_in[9]),
        .I3(\r_reg[iforce][0]__0 [8]),
        .I4(p_5_in[9]),
        .I5(\r_reg[imask][0]__0 [8]),
        .O(\r[irl][0][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_5 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][0]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][0]__0 [7]),
        .O(\r[irl][0][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \r[irl][0][3]_i_6 
       (.I0(\r[irl][0][3]_i_15_n_0 ),
        .I1(\r[irl][0][3]_i_16_n_0 ),
        .I2(\r[irl][0][2]_i_7_n_0 ),
        .I3(\r[irl][0][2]_i_8_n_0 ),
        .I4(\r[irl][0][2]_i_9_n_0 ),
        .I5(\r[irl][0][2]_i_10_n_0 ),
        .O(\r[irl][0][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_7 
       (.I0(p_6_in[1]),
        .I1(\r_reg[iforce][0]__0 [0]),
        .I2(p_5_in[1]),
        .I3(\r_reg[imask][0]__0 [0]),
        .O(\r[irl][0][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_8 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][0]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][0]__0 [2]),
        .O(\r[irl][0][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][0][3]_i_9 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][0]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][0]__0 [3]),
        .O(\r[irl][0][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCCAAC0AA)) 
    \r[irl][1][0]_i_1 
       (.I0(\r[irl][1][0]_i_2_n_0 ),
        .I1(\r[irl][1][0]_i_3_n_0 ),
        .I2(\r[irl][1][0]_i_4_n_0 ),
        .I3(\r[irl][1][3]_i_3_n_0 ),
        .I4(\r[irl][1][3]_i_4_n_0 ),
        .O(\r[irl][1][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF007500FF)) 
    \r[irl][1][0]_i_2 
       (.I0(\r[irl][1][1]_i_4_n_0 ),
        .I1(\r[irl][1][3]_i_10_n_0 ),
        .I2(p_6_in[3]),
        .I3(\r[irl][1][0]_i_5_n_0 ),
        .I4(\r[irl][1][3]_i_8_n_0 ),
        .I5(\r[irl][1][3]_i_9_n_0 ),
        .O(\r[irl][1][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEEF)) 
    \r[irl][1][0]_i_3 
       (.I0(\r[irl][1][3]_i_5_n_0 ),
        .I1(\r[irl][1][1]_i_8_n_0 ),
        .I2(p_6_in[1]),
        .I3(\r[irl][1][0]_i_6_n_0 ),
        .I4(\r[irl][1][3]_i_11_n_0 ),
        .I5(\r[irl][1][2]_i_18_n_0 ),
        .O(\r[irl][1][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5400FFFF54000000)) 
    \r[irl][1][0]_i_4 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][1]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][1]__0 [2]),
        .I4(\r[irl][1][2]_i_5_n_0 ),
        .I5(\r[irl][1][0]_i_7_n_0 ),
        .O(\r[irl][1][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0FFF0F0F0F2)) 
    \r[irl][1][0]_i_5 
       (.I0(\r[irl][1][2]_i_11_n_0 ),
        .I1(\r[irl][1][3]_i_18_n_0 ),
        .I2(\r[irl][1][0]_i_8_n_0 ),
        .I3(\r[irl][1][3]_i_17_n_0 ),
        .I4(\r[irl][1][3]_i_7_n_0 ),
        .I5(\r[irl][1][3]_i_6_n_0 ),
        .O(\r[irl][1][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][0]_i_6 
       (.I0(\r_reg[imask][1]__0 [0]),
        .I1(p_5_in[1]),
        .I2(\r_reg[iforce][1]__0 [0]),
        .O(\r[irl][1][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEF0F0FFF0F0F0)) 
    \r[irl][1][0]_i_7 
       (.I0(\r[irl][1][0]_i_9_n_0 ),
        .I1(\r[irl][1][3]_i_20_n_0 ),
        .I2(\r[irl][1][2]_i_13_n_0 ),
        .I3(\r[irl][1][2]_i_15_n_0 ),
        .I4(\r[irl][1][2]_i_14_n_0 ),
        .I5(\r[irl][1][1]_i_16_n_0 ),
        .O(\r[irl][1][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF000FC00F000FE00)) 
    \r[irl][1][0]_i_8 
       (.I0(\r[irl][1][3]_i_14_n_0 ),
        .I1(\r[irl][1][2]_i_9_n_0 ),
        .I2(\r[irl][1][2]_i_8_n_0 ),
        .I3(\r[irl][1][2]_i_7_n_0 ),
        .I4(\r[irl][1][3]_i_16_n_0 ),
        .I5(\r[irl][1][3]_i_15_n_0 ),
        .O(\r[irl][1][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88888A888A8A8A8A)) 
    \r[irl][1][0]_i_9 
       (.I0(\r[irl][1][3]_i_19_n_0 ),
        .I1(\r[irl][1][2]_i_17_n_0 ),
        .I2(\r[irl][1][3]_i_12_n_0 ),
        .I3(\r[irl][1][2]_i_20_n_0 ),
        .I4(\r[irl][1][2]_i_21_n_0 ),
        .I5(\r[irl][1][2]_i_22_n_0 ),
        .O(\r[irl][1][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAFFAAF0AAFFAAF3)) 
    \r[irl][1][1]_i_1 
       (.I0(\r[irl][1][1]_i_2_n_0 ),
        .I1(\r[irl][1][1]_i_3_n_0 ),
        .I2(\r[irl][1][1]_i_4_n_0 ),
        .I3(\r[irl][1][2]_i_3_n_0 ),
        .I4(\r[irl][1][1]_i_5_n_0 ),
        .I5(\r[irl][1][1]_i_6_n_0 ),
        .O(\r[irl][1][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00A8FFFF)) 
    \r[irl][1][1]_i_10 
       (.I0(\r_reg[imask][1]__0 [8]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][1]__0 [8]),
        .I3(p_6_in[9]),
        .I4(\r[irl][1][3]_i_13_n_0 ),
        .O(\r[irl][1][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F000F0E0F000F0)) 
    \r[irl][1][1]_i_11 
       (.I0(\r[irl][1][2]_i_17_n_0 ),
        .I1(\r[irl][1][3]_i_12_n_0 ),
        .I2(\r[irl][1][1]_i_15_n_0 ),
        .I3(\r[irl][1][1]_i_16_n_0 ),
        .I4(\r[irl][1][3]_i_19_n_0 ),
        .I5(\r[irl][1][3]_i_20_n_0 ),
        .O(\r[irl][1][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][1]_i_12 
       (.I0(\r_reg[imask][1]__0 [10]),
        .I1(p_5_in[11]),
        .I2(\r_reg[iforce][1]__0 [10]),
        .O(\r[irl][1][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000777F)) 
    \r[irl][1][1]_i_13 
       (.I0(p_6_in[15]),
        .I1(\r_reg[imask][1]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[iforce][1]__0 [14]),
        .I4(\r[irl][1][2]_i_8_n_0 ),
        .O(\r[irl][1][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][1][1]_i_14 
       (.I0(\r_reg[imask][1]__0 [6]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][1]__0 [6]),
        .I3(p_6_in[7]),
        .I4(\r[irl][1][2]_i_21_n_0 ),
        .O(\r[irl][1][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][1][1]_i_15 
       (.I0(\r_reg[imask][1]__0 [13]),
        .I1(p_5_in[14]),
        .I2(\r_reg[iforce][1]__0 [13]),
        .I3(p_6_in[14]),
        .I4(\r[irl][1][2]_i_13_n_0 ),
        .O(\r[irl][1][1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][1][1]_i_16 
       (.I0(\r_reg[imask][1]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][1]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][1][2]_i_15_n_0 ),
        .O(\r[irl][1][1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00F4F4)) 
    \r[irl][1][1]_i_2 
       (.I0(\r[irl][1][2]_i_12_n_0 ),
        .I1(p_6_in[7]),
        .I2(\r[irl][1][2]_i_11_n_0 ),
        .I3(\r[irl][1][1]_i_7_n_0 ),
        .I4(\r[irl][1][3]_i_2_n_0 ),
        .O(\r[irl][1][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF1111000F)) 
    \r[irl][1][1]_i_3 
       (.I0(\r[irl][1][1]_i_8_n_0 ),
        .I1(\r[irl][1][3]_i_11_n_0 ),
        .I2(\r[irl][1][1]_i_9_n_0 ),
        .I3(\r[irl][1][1]_i_10_n_0 ),
        .I4(\r[irl][1][2]_i_5_n_0 ),
        .I5(\r[irl][1][1]_i_11_n_0 ),
        .O(\r[irl][1][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][1]_i_4 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][1]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][1]__0 [1]),
        .O(\r[irl][1][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][1]_i_5 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][1]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][1]__0 [2]),
        .O(\r[irl][1][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][1]_i_6 
       (.I0(p_6_in[1]),
        .I1(\r_reg[iforce][1]__0 [0]),
        .I2(p_5_in[1]),
        .I3(\r_reg[imask][1]__0 [0]),
        .O(\r[irl][1][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF400F4FF)) 
    \r[irl][1][1]_i_7 
       (.I0(\r[irl][1][1]_i_12_n_0 ),
        .I1(p_6_in[11]),
        .I2(\r[irl][1][3]_i_14_n_0 ),
        .I3(\r[irl][1][2]_i_2_n_0 ),
        .I4(\r[irl][1][1]_i_13_n_0 ),
        .O(\r[irl][1][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][1]_i_8 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][1]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][1]__0 [1]),
        .O(\r[irl][1][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][1][1]_i_9 
       (.I0(\r_reg[imask][1]__0 [7]),
        .I1(p_5_in[8]),
        .I2(\r_reg[iforce][1]__0 [7]),
        .I3(p_6_in[8]),
        .I4(\r[irl][1][1]_i_14_n_0 ),
        .O(\r[irl][1][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7070707070FF7070)) 
    \r[irl][1][2]_i_1 
       (.I0(\r[irl][1][2]_i_2_n_0 ),
        .I1(\r[irl][1][3]_i_2_n_0 ),
        .I2(\r[irl][1][2]_i_3_n_0 ),
        .I3(\r[irl][1][2]_i_4_n_0 ),
        .I4(\r[irl][1][3]_i_3_n_0 ),
        .I5(\r[irl][1][2]_i_5_n_0 ),
        .O(\r[irl][1][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][2]_i_10 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][1]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][1]__0 [4]),
        .O(\r[irl][1][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][2]_i_11 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][1]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][1]__0 [5]),
        .O(\r[irl][1][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][2]_i_12 
       (.I0(\r_reg[imask][1]__0 [6]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][1]__0 [6]),
        .O(\r[irl][1][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][2]_i_13 
       (.I0(p_6_in[15]),
        .I1(\r_reg[iforce][1]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[imask][1]__0 [14]),
        .O(\r[irl][1][2]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFF)) 
    \r[irl][1][2]_i_14 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][1]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][1]__0 [13]),
        .O(\r[irl][1][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][2]_i_15 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][1]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][1]__0 [12]),
        .O(\r[irl][1][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][2]_i_16 
       (.I0(\r_reg[imask][1]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][1]__0 [11]),
        .O(\r[irl][1][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][2]_i_17 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][1]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][1]__0 [8]),
        .O(\r[irl][1][2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF1FFFF)) 
    \r[irl][1][2]_i_18 
       (.I0(p_6_in[4]),
        .I1(\r[irl][1][2]_i_19_n_0 ),
        .I2(\r[irl][1][2]_i_20_n_0 ),
        .I3(\r[irl][1][2]_i_21_n_0 ),
        .I4(\r[irl][1][2]_i_22_n_0 ),
        .O(\r[irl][1][2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][2]_i_19 
       (.I0(\r_reg[imask][1]__0 [3]),
        .I1(p_5_in[4]),
        .I2(\r_reg[iforce][1]__0 [3]),
        .O(\r[irl][1][2]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000000D0)) 
    \r[irl][1][2]_i_2 
       (.I0(p_6_in[13]),
        .I1(\r[irl][1][2]_i_6_n_0 ),
        .I2(\r[irl][1][2]_i_7_n_0 ),
        .I3(\r[irl][1][2]_i_8_n_0 ),
        .I4(\r[irl][1][2]_i_9_n_0 ),
        .O(\r[irl][1][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][2]_i_20 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][1]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][1]__0 [4]),
        .O(\r[irl][1][2]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][2]_i_21 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][1]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][1]__0 [5]),
        .O(\r[irl][1][2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFF)) 
    \r[irl][1][2]_i_22 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][1]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][1]__0 [6]),
        .O(\r[irl][1][2]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000001010001))
    \r[irl][1][2]_i_3 
       (.I0(\r[irl][1][3]_i_9_n_0 ),
        .I1(\r[irl][1][2]_i_10_n_0 ),
        .I2(\r[irl][1][2]_i_11_n_0 ),
        .I3(p_6_in[7]),
        .I4(\r[irl][1][2]_i_12_n_0 ),
        .I5(\r[irl][1][3]_i_2_n_0 ),
        .O(\r[irl][1][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0404040000000000)) 
    \r[irl][1][2]_i_4 
       (.I0(\r[irl][1][2]_i_13_n_0 ),
        .I1(\r[irl][1][2]_i_14_n_0 ),
        .I2(\r[irl][1][2]_i_15_n_0 ),
        .I3(p_6_in[12]),
        .I4(\r[irl][1][2]_i_16_n_0 ),
        .I5(\r[irl][1][3]_i_5_n_0 ),
        .O(\r[irl][1][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \r[irl][1][2]_i_5 
       (.I0(\r[irl][1][2]_i_17_n_0 ),
        .I1(\r[irl][1][3]_i_13_n_0 ),
        .I2(\r[irl][1][3]_i_12_n_0 ),
        .I3(\r[irl][1][2]_i_18_n_0 ),
        .O(\r[irl][1][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][2]_i_6 
       (.I0(\r_reg[imask][1]__0 [12]),
        .I1(p_5_in[13]),
        .I2(\r_reg[iforce][1]__0 [12]),
        .O(\r[irl][1][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1FFF)) 
    \r[irl][1][2]_i_7 
       (.I0(\r_reg[iforce][1]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[imask][1]__0 [14]),
        .I3(p_6_in[15]),
        .O(\r[irl][1][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][2]_i_8 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][1]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][1]__0 [13]),
        .O(\r[irl][1][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][2]_i_9 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][1]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][1]__0 [11]),
        .O(\r[irl][1][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hAEAA)) 
    \r[irl][1][3]_i_1 
       (.I0(\r[irl][1][3]_i_2_n_0 ),
        .I1(\r[irl][1][3]_i_3_n_0 ),
        .I2(\r[irl][1][3]_i_4_n_0 ),
        .I3(\r[irl][1][3]_i_5_n_0 ),
        .O(\r[irl][1][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][1][3]_i_10 
       (.I0(\r_reg[imask][1]__0 [2]),
        .I1(p_5_in[3]),
        .I2(\r_reg[iforce][1]__0 [2]),
        .O(\r[irl][1][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][3]_i_11 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][1]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][1]__0 [2]),
        .O(\r[irl][1][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][3]_i_12 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][1]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][1]__0 [7]),
        .O(\r[irl][1][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \r[irl][1][3]_i_13 
       (.I0(\r[irl][1][3]_i_19_n_0 ),
        .I1(\r[irl][1][3]_i_20_n_0 ),
        .I2(\r[irl][1][2]_i_13_n_0 ),
        .I3(\r[irl][1][2]_i_14_n_0 ),
        .I4(\r[irl][1][2]_i_15_n_0 ),
        .I5(\r[irl][1][3]_i_21_n_0 ),
        .O(\r[irl][1][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_14 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][1]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][1]__0 [9]),
        .O(\r[irl][1][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_15 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][1]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][1]__0 [10]),
        .O(\r[irl][1][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_16 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][1]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][1]__0 [12]),
        .O(\r[irl][1][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_17 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][1]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][1]__0 [8]),
        .O(\r[irl][1][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_18 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][1]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][1]__0 [6]),
        .O(\r[irl][1][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFF)) 
    \r[irl][1][3]_i_19 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][1]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][1]__0 [9]),
        .O(\r[irl][1][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][1][3]_i_2 
       (.I0(\r[irl][1][3]_i_6_n_0 ),
        .I1(p_6_in[9]),
        .I2(\r_reg[iforce][1]__0 [8]),
        .I3(p_5_in[9]),
        .I4(\r_reg[imask][1]__0 [8]),
        .I5(\r[irl][1][3]_i_7_n_0 ),
        .O(\r[irl][1][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][3]_i_20 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][1]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][1]__0 [10]),
        .O(\r[irl][1][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][1][3]_i_21 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][1]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][1]__0 [11]),
        .O(\r[irl][1][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000004000404)) 
    \r[irl][1][3]_i_3 
       (.I0(\r[irl][1][1]_i_4_n_0 ),
        .I1(\r[irl][1][3]_i_8_n_0 ),
        .I2(\r[irl][1][3]_i_9_n_0 ),
        .I3(\r[irl][1][3]_i_10_n_0 ),
        .I4(p_6_in[3]),
        .I5(\r[irl][1][1]_i_6_n_0 ),
        .O(\r[irl][1][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444404040444)) 
    \r[irl][1][3]_i_4 
       (.I0(\r[irl][1][3]_i_11_n_0 ),
        .I1(\r[irl][1][2]_i_5_n_0 ),
        .I2(\r_reg[imask][1]__0 [1]),
        .I3(p_5_in[2]),
        .I4(\r_reg[iforce][1]__0 [1]),
        .I5(p_6_in[2]),
        .O(\r[irl][1][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFBFBFBBBBBBBBBB)) 
    \r[irl][1][3]_i_5 
       (.I0(\r[irl][1][3]_i_12_n_0 ),
        .I1(\r[irl][1][3]_i_13_n_0 ),
        .I2(p_6_in[9]),
        .I3(\r_reg[iforce][1]__0 [8]),
        .I4(p_5_in[9]),
        .I5(\r_reg[imask][1]__0 [8]),
        .O(\r[irl][1][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_6 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][1]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][1]__0 [7]),
        .O(\r[irl][1][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \r[irl][1][3]_i_7 
       (.I0(\r[irl][1][3]_i_14_n_0 ),
        .I1(\r[irl][1][3]_i_15_n_0 ),
        .I2(\r[irl][1][3]_i_16_n_0 ),
        .I3(\r[irl][1][2]_i_7_n_0 ),
        .I4(\r[irl][1][2]_i_8_n_0 ),
        .I5(\r[irl][1][2]_i_9_n_0 ),
        .O(\r[irl][1][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[irl][1][3]_i_8 
       (.I0(\r[irl][1][3]_i_7_n_0 ),
        .I1(\r[irl][1][3]_i_17_n_0 ),
        .I2(\r[irl][1][3]_i_6_n_0 ),
        .I3(\r[irl][1][3]_i_18_n_0 ),
        .I4(\r[irl][1][2]_i_11_n_0 ),
        .I5(\r[irl][1][2]_i_10_n_0 ),
        .O(\r[irl][1][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][1][3]_i_9 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][1]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][1]__0 [3]),
        .O(\r[irl][1][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF1B1B00FF)) 
    \r[irl][2][0]_i_1 
       (.I0(\r[irl][2][1]_i_6_n_0 ),
        .I1(\r[irl][2][1]_i_7_n_0 ),
        .I2(\r[irl][2][0]_i_2_n_0 ),
        .I3(\r[irl][2][0]_i_3_n_0 ),
        .I4(\r[irl][2][3]_i_4_n_0 ),
        .I5(\r[irl][2][0]_i_4_n_0 ),
        .O(\r[irl][2][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][2][0]_i_10 
       (.I0(\r_reg[imask][2]__0 [10]),
        .I1(p_5_in[11]),
        .I2(\r_reg[iforce][2]__0 [10]),
        .O(\r[irl][2][0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF000000FF00BA00)) 
    \r[irl][2][0]_i_11 
       (.I0(\r[irl][2][2]_i_9_n_0 ),
        .I1(\r[irl][2][3]_i_17_n_0 ),
        .I2(\r[irl][2][0]_i_13_n_0 ),
        .I3(\r[irl][2][2]_i_8_n_0 ),
        .I4(\r[irl][2][2]_i_7_n_0 ),
        .I5(\r[irl][2][0]_i_14_n_0 ),
        .O(\r[irl][2][0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \r[irl][2][0]_i_12 
       (.I0(\r[irl][2][2]_i_9_n_0 ),
        .I1(\r[irl][2][2]_i_8_n_0 ),
        .I2(\r[irl][2][2]_i_7_n_0 ),
        .I3(\r[irl][2][0]_i_14_n_0 ),
        .I4(\r[irl][2][3]_i_17_n_0 ),
        .I5(\r[irl][2][0]_i_13_n_0 ),
        .O(\r[irl][2][0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][0]_i_13 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][2]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][2]__0 [9]),
        .O(\r[irl][2][0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][0]_i_14 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][2]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][2]__0 [12]),
        .O(\r[irl][2][0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8888B888B8B8B8B8)) 
    \r[irl][2][0]_i_2 
       (.I0(\r[irl][2][1]_i_15_n_0 ),
        .I1(\r[irl][2][2]_i_11_n_0 ),
        .I2(\r[irl][2][0]_i_5_n_0 ),
        .I3(\r[irl][2][0]_i_6_n_0 ),
        .I4(\r[irl][2][0]_i_7_n_0 ),
        .I5(\r[irl][2][3]_i_3_n_0 ),
        .O(\r[irl][2][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0FFF0F0F0F4)) 
    \r[irl][2][0]_i_3 
       (.I0(\r[irl][2][3]_i_16_n_0 ),
        .I1(\r[irl][2][3]_i_12_n_0 ),
        .I2(\r[irl][2][0]_i_8_n_0 ),
        .I3(\r[irl][2][3]_i_14_n_0 ),
        .I4(\r[irl][2][3]_i_13_n_0 ),
        .I5(\r[irl][2][3]_i_15_n_0 ),
        .O(\r[irl][2][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0002)) 
    \r[irl][2][0]_i_4 
       (.I0(\r[irl][2][1]_i_14_n_0 ),
        .I1(\r[irl][2][1]_i_12_n_0 ),
        .I2(\r[irl][2][1]_i_13_n_0 ),
        .I3(\r[irl][2][1]_i_11_n_0 ),
        .O(\r[irl][2][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7774444477747774)) 
    \r[irl][2][0]_i_5 
       (.I0(\r[irl][2][0]_i_9_n_0 ),
        .I1(\r[irl][2][2]_i_10_n_0 ),
        .I2(\r[irl][2][0]_i_10_n_0 ),
        .I3(p_6_in[11]),
        .I4(\r[irl][2][3]_i_9_n_0 ),
        .I5(\r[irl][2][3]_i_10_n_0 ),
        .O(\r[irl][2][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][0]_i_6 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][2]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][2]__0 [5]),
        .O(\r[irl][2][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][0]_i_7 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][2]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][2]__0 [6]),
        .O(\r[irl][2][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0FFF0F0F0F2F0F0)) 
    \r[irl][2][0]_i_8 
       (.I0(\r[irl][2][1]_i_9_n_0 ),
        .I1(\r[irl][2][1]_i_10_n_0 ),
        .I2(\r[irl][2][0]_i_11_n_0 ),
        .I3(\r[irl][2][3]_i_23_n_0 ),
        .I4(\r[irl][2][0]_i_12_n_0 ),
        .I5(\r[irl][2][3]_i_5_n_0 ),
        .O(\r[irl][2][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF00A800A800A8)) 
    \r[irl][2][0]_i_9 
       (.I0(\r_reg[imask][2]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[iforce][2]__0 [14]),
        .I3(p_6_in[15]),
        .I4(\r[irl][2][3]_i_19_n_0 ),
        .I5(\r[irl][2][3]_i_21_n_0 ),
        .O(\r[irl][2][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5503550355035500)) 
    \r[irl][2][1]_i_1 
       (.I0(\r[irl][2][1]_i_2_n_0 ),
        .I1(\r[irl][2][1]_i_3_n_0 ),
        .I2(\r[irl][2][1]_i_4_n_0 ),
        .I3(\r[irl][2][1]_i_5_n_0 ),
        .I4(\r[irl][2][1]_i_6_n_0 ),
        .I5(\r[irl][2][1]_i_7_n_0 ),
        .O(\r[irl][2][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][1]_i_10 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][2]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][2]__0 [6]),
        .O(\r[irl][2][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][1]_i_11 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][2]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][2]__0 [2]),
        .O(\r[irl][2][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEEFEFEFEEE)) 
    \r[irl][2][1]_i_12 
       (.I0(\r[irl][2][1]_i_7_n_0 ),
        .I1(\r[irl][2][1]_i_15_n_0 ),
        .I2(\r_reg[imask][2]__0 [0]),
        .I3(p_5_in[1]),
        .I4(\r_reg[iforce][2]__0 [0]),
        .I5(p_6_in[1]),
        .O(\r[irl][2][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][1]_i_13 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][2]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][2]__0 [4]),
        .O(\r[irl][2][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    \r[irl][2][1]_i_14 
       (.I0(\r[irl][2][3]_i_11_n_0 ),
        .I1(\r[irl][2][3]_i_10_n_0 ),
        .I2(\r[irl][2][3]_i_9_n_0 ),
        .I3(\r[irl][2][2]_i_12_n_0 ),
        .I4(\r[irl][2][3]_i_8_n_0 ),
        .O(\r[irl][2][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][1]_i_15 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][2]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][2]__0 [3]),
        .O(\r[irl][2][1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0303030F0303030B)) 
    \r[irl][2][1]_i_16 
       (.I0(\r[irl][2][2]_i_12_n_0 ),
        .I1(\r[irl][2][1]_i_19_n_0 ),
        .I2(\r[irl][2][1]_i_20_n_0 ),
        .I3(\r[irl][2][3]_i_22_n_0 ),
        .I4(\r[irl][2][3]_i_9_n_0 ),
        .I5(\r[irl][2][1]_i_21_n_0 ),
        .O(\r[irl][2][1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][2][1]_i_17 
       (.I0(\r_reg[imask][2]__0 [4]),
        .I1(p_5_in[5]),
        .I2(\r_reg[iforce][2]__0 [4]),
        .O(\r[irl][2][1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA800FFFF)) 
    \r[irl][2][1]_i_18 
       (.I0(\r_reg[imask][2]__0 [13]),
        .I1(p_5_in[14]),
        .I2(\r_reg[iforce][2]__0 [13]),
        .I3(p_6_in[14]),
        .I4(\r[irl][2][2]_i_8_n_0 ),
        .O(\r[irl][2][1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][2][1]_i_19 
       (.I0(\r_reg[imask][2]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][2]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][2][3]_i_19_n_0 ),
        .O(\r[irl][2][1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00F000F000F00EFE)) 
    \r[irl][2][1]_i_2 
       (.I0(\r[irl][2][3]_i_14_n_0 ),
        .I1(\r[irl][2][3]_i_15_n_0 ),
        .I2(\r[irl][2][3]_i_2_n_0 ),
        .I3(\r[irl][2][1]_i_8_n_0 ),
        .I4(\r[irl][2][1]_i_9_n_0 ),
        .I5(\r[irl][2][1]_i_10_n_0 ),
        .O(\r[irl][2][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00A8FFFF)) 
    \r[irl][2][1]_i_20 
       (.I0(\r_reg[imask][2]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[iforce][2]__0 [14]),
        .I3(p_6_in[15]),
        .I4(\r[irl][2][3]_i_21_n_0 ),
        .O(\r[irl][2][1]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00A8)) 
    \r[irl][2][1]_i_21 
       (.I0(\r_reg[imask][2]__0 [7]),
        .I1(p_5_in[8]),
        .I2(\r_reg[iforce][2]__0 [7]),
        .I3(p_6_in[8]),
        .I4(\r[irl][2][3]_i_10_n_0 ),
        .O(\r[irl][2][1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF1FF01000100)) 
    \r[irl][2][1]_i_3 
       (.I0(\r[irl][2][1]_i_11_n_0 ),
        .I1(\r[irl][2][1]_i_12_n_0 ),
        .I2(\r[irl][2][1]_i_13_n_0 ),
        .I3(\r[irl][2][1]_i_14_n_0 ),
        .I4(\r[irl][2][1]_i_15_n_0 ),
        .I5(\r[irl][2][1]_i_16_n_0 ),
        .O(\r[irl][2][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][1]_i_4 
       (.I0(p_6_in[1]),
        .I1(\r_reg[iforce][2]__0 [0]),
        .I2(p_5_in[1]),
        .I3(\r_reg[imask][2]__0 [0]),
        .O(\r[irl][2][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFEEFE)) 
    \r[irl][2][1]_i_5 
       (.I0(\r[irl][2][3]_i_16_n_0 ),
        .I1(\r[irl][2][3]_i_15_n_0 ),
        .I2(p_6_in[5]),
        .I3(\r[irl][2][1]_i_17_n_0 ),
        .I4(\r[irl][2][3]_i_13_n_0 ),
        .I5(\r[irl][2][3]_i_12_n_0 ),
        .O(\r[irl][2][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF00A8FFFFFFFF)) 
    \r[irl][2][1]_i_6 
       (.I0(\r_reg[imask][2]__0 [2]),
        .I1(p_5_in[3]),
        .I2(\r_reg[iforce][2]__0 [2]),
        .I3(p_6_in[3]),
        .I4(\r[irl][2][1]_i_15_n_0 ),
        .I5(\r[irl][2][2]_i_11_n_0 ),
        .O(\r[irl][2][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][1]_i_7 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][2]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][2]__0 [1]),
        .O(\r[irl][2][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r[irl][2][1]_i_8 
       (.I0(\r[irl][2][3]_i_7_n_0 ),
        .I1(\r[irl][2][2]_i_2_n_0 ),
        .I2(\r[irl][2][1]_i_18_n_0 ),
        .O(\r[irl][2][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][1]_i_9 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][2]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][2]__0 [5]),
        .O(\r[irl][2][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7070707070FF7070)) 
    \r[irl][2][2]_i_1 
       (.I0(\r[irl][2][2]_i_2_n_0 ),
        .I1(\r[irl][2][3]_i_2_n_0 ),
        .I2(\r[irl][2][2]_i_3_n_0 ),
        .I3(\r[irl][2][2]_i_4_n_0 ),
        .I4(\r[irl][2][3]_i_4_n_0 ),
        .I5(\r[irl][2][2]_i_5_n_0 ),
        .O(\r[irl][2][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFDFDFDFF)) 
    \r[irl][2][2]_i_10 
       (.I0(\r[irl][2][3]_i_21_n_0 ),
        .I1(\r[irl][2][3]_i_20_n_0 ),
        .I2(\r[irl][2][3]_i_19_n_0 ),
        .I3(p_6_in[12]),
        .I4(\r[irl][2][3]_i_18_n_0 ),
        .O(\r[irl][2][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \r[irl][2][2]_i_11 
       (.I0(\r[irl][2][3]_i_8_n_0 ),
        .I1(\r[irl][2][2]_i_12_n_0 ),
        .I2(\r[irl][2][3]_i_9_n_0 ),
        .I3(\r[irl][2][3]_i_10_n_0 ),
        .I4(\r[irl][2][3]_i_11_n_0 ),
        .I5(\r[irl][2][1]_i_13_n_0 ),
        .O(\r[irl][2][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][2][2]_i_12 
       (.I0(\r_reg[imask][2]__0 [6]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][2]__0 [6]),
        .I3(p_6_in[7]),
        .I4(\r[irl][2][0]_i_6_n_0 ),
        .O(\r[irl][2][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000D00)) 
    \r[irl][2][2]_i_2 
       (.I0(p_6_in[13]),
        .I1(\r[irl][2][2]_i_6_n_0 ),
        .I2(\r[irl][2][2]_i_7_n_0 ),
        .I3(\r[irl][2][2]_i_8_n_0 ),
        .I4(\r[irl][2][2]_i_9_n_0 ),
        .O(\r[irl][2][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][2][2]_i_3 
       (.I0(\r[irl][2][3]_i_15_n_0 ),
        .I1(p_6_in[5]),
        .I2(\r_reg[iforce][2]__0 [4]),
        .I3(p_5_in[5]),
        .I4(\r_reg[imask][2]__0 [4]),
        .I5(\r[irl][2][3]_i_13_n_0 ),
        .O(\r[irl][2][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \r[irl][2][2]_i_4 
       (.I0(\r[irl][2][2]_i_10_n_0 ),
        .I1(\r[irl][2][3]_i_3_n_0 ),
        .O(\r[irl][2][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAA222A)) 
    \r[irl][2][2]_i_5 
       (.I0(\r[irl][2][2]_i_11_n_0 ),
        .I1(\r_reg[imask][2]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[iforce][2]__0 [3]),
        .I4(p_6_in[4]),
        .O(\r[irl][2][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][2][2]_i_6 
       (.I0(\r_reg[imask][2]__0 [12]),
        .I1(p_5_in[13]),
        .I2(\r_reg[iforce][2]__0 [12]),
        .O(\r[irl][2][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][2]_i_7 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][2]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][2]__0 [13]),
        .O(\r[irl][2][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1FFF)) 
    \r[irl][2][2]_i_8 
       (.I0(\r_reg[iforce][2]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[imask][2]__0 [14]),
        .I3(p_6_in[15]),
        .O(\r[irl][2][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][2]_i_9 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][2]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][2]__0 [11]),
        .O(\r[irl][2][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    \r[irl][2][3]_i_1 
       (.I0(\r[irl][2][3]_i_2_n_0 ),
        .I1(\r[irl][2][3]_i_3_n_0 ),
        .I2(\r[irl][2][3]_i_4_n_0 ),
        .O(\r[irl][2][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_10 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][2]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][2]__0 [8]),
        .O(\r[irl][2][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_11 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][2]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][2]__0 [7]),
        .O(\r[irl][2][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_12 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][2]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][2]__0 [1]),
        .O(\r[irl][2][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFEFFFF)) 
    \r[irl][2][3]_i_13 
       (.I0(\r[irl][2][1]_i_9_n_0 ),
        .I1(\r[irl][2][1]_i_10_n_0 ),
        .I2(\r[irl][2][3]_i_5_n_0 ),
        .I3(\r[irl][2][3]_i_23_n_0 ),
        .I4(\r[irl][2][2]_i_2_n_0 ),
        .I5(\r[irl][2][3]_i_7_n_0 ),
        .O(\r[irl][2][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_14 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][2]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][2]__0 [4]),
        .O(\r[irl][2][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_15 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][2]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][2]__0 [3]),
        .O(\r[irl][2][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_16 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][2]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][2]__0 [2]),
        .O(\r[irl][2][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_17 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][2]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][2]__0 [10]),
        .O(\r[irl][2][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][2][3]_i_18 
       (.I0(\r_reg[imask][2]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][2]__0 [11]),
        .O(\r[irl][2][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_19 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][2]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][2]__0 [12]),
        .O(\r[irl][2][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFAEFF)) 
    \r[irl][2][3]_i_2 
       (.I0(\r[irl][2][3]_i_5_n_0 ),
        .I1(p_6_in[9]),
        .I2(\r[irl][2][3]_i_6_n_0 ),
        .I3(\r[irl][2][2]_i_2_n_0 ),
        .I4(\r[irl][2][3]_i_7_n_0 ),
        .O(\r[irl][2][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_20 
       (.I0(p_6_in[15]),
        .I1(\r_reg[iforce][2]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[imask][2]__0 [14]),
        .O(\r[irl][2][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFF)) 
    \r[irl][2][3]_i_21 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][2]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][2]__0 [13]),
        .O(\r[irl][2][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_22 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][2]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][2]__0 [10]),
        .O(\r[irl][2][3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_23 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][2]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][2]__0 [8]),
        .O(\r[irl][2][3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[irl][2][3]_i_3 
       (.I0(\r[irl][2][3]_i_8_n_0 ),
        .I1(\r[irl][2][3]_i_9_n_0 ),
        .I2(\r[irl][2][3]_i_10_n_0 ),
        .I3(\r[irl][2][3]_i_11_n_0 ),
        .O(\r[irl][2][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[irl][2][3]_i_4 
       (.I0(\r[irl][2][3]_i_12_n_0 ),
        .I1(\r[irl][2][3]_i_13_n_0 ),
        .I2(\r[irl][2][3]_i_14_n_0 ),
        .I3(\r[irl][2][3]_i_15_n_0 ),
        .I4(\r[irl][2][3]_i_16_n_0 ),
        .I5(\r[irl][2][1]_i_4_n_0 ),
        .O(\r[irl][2][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][2][3]_i_5 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][2]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][2]__0 [7]),
        .O(\r[irl][2][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][2][3]_i_6 
       (.I0(\r_reg[imask][2]__0 [8]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][2]__0 [8]),
        .O(\r[irl][2][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA800)) 
    \r[irl][2][3]_i_7 
       (.I0(\r_reg[imask][2]__0 [9]),
        .I1(p_5_in[10]),
        .I2(\r_reg[iforce][2]__0 [9]),
        .I3(p_6_in[10]),
        .I4(\r[irl][2][3]_i_17_n_0 ),
        .O(\r[irl][2][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF1FFFF)) 
    \r[irl][2][3]_i_8 
       (.I0(\r[irl][2][3]_i_18_n_0 ),
        .I1(p_6_in[12]),
        .I2(\r[irl][2][3]_i_19_n_0 ),
        .I3(\r[irl][2][3]_i_20_n_0 ),
        .I4(\r[irl][2][3]_i_21_n_0 ),
        .I5(\r[irl][2][3]_i_22_n_0 ),
        .O(\r[irl][2][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][2][3]_i_9 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][2]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][2]__0 [9]),
        .O(\r[irl][2][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0303AAAAFF00AAAA)) 
    \r[irl][3][0]_i_1 
       (.I0(\r[irl][3][0]_i_2_n_0 ),
        .I1(p_6_in[1]),
        .I2(\r[irl][3][0]_i_3_n_0 ),
        .I3(\r[irl][3][0]_i_4_n_0 ),
        .I4(\r[irl][3][3]_i_3_n_0 ),
        .I5(\r[irl][3][1]_i_6_n_0 ),
        .O(\r[irl][3][0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF004F00FF)) 
    \r[irl][3][0]_i_2 
       (.I0(\r[irl][3][3]_i_10_n_0 ),
        .I1(p_6_in[3]),
        .I2(\r[irl][3][3]_i_7_n_0 ),
        .I3(\r[irl][3][0]_i_5_n_0 ),
        .I4(\r[irl][3][3]_i_8_n_0 ),
        .I5(\r[irl][3][3]_i_9_n_0 ),
        .O(\r[irl][3][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][0]_i_3 
       (.I0(\r_reg[imask][3]__0 [0]),
        .I1(p_5_in[1]),
        .I2(\r_reg[iforce][3]__0 [0]),
        .O(\r[irl][3][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00C000E00FCF0FEF)) 
    \r[irl][3][0]_i_4 
       (.I0(\r[irl][3][1]_i_13_n_0 ),
        .I1(\r[irl][3][2]_i_13_n_0 ),
        .I2(\r[irl][3][0]_i_6_n_0 ),
        .I3(\r[irl][3][2]_i_16_n_0 ),
        .I4(\r[irl][3][2]_i_17_n_0 ),
        .I5(\r[irl][3][0]_i_7_n_0 ),
        .O(\r[irl][3][0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF0F0F0FFF0F0F0F2)) 
    \r[irl][3][0]_i_5 
       (.I0(\r[irl][3][1]_i_8_n_0 ),
        .I1(\r[irl][3][3]_i_16_n_0 ),
        .I2(\r[irl][3][0]_i_8_n_0 ),
        .I3(\r[irl][3][3]_i_15_n_0 ),
        .I4(\r[irl][3][3]_i_6_n_0 ),
        .I5(\r[irl][3][3]_i_5_n_0 ),
        .O(\r[irl][3][0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000E000E000E0000)) 
    \r[irl][3][0]_i_6 
       (.I0(p_6_in[7]),
        .I1(\r[irl][3][1]_i_7_n_0 ),
        .I2(\r[irl][3][3]_i_11_n_0 ),
        .I3(\r[irl][3][3]_i_12_n_0 ),
        .I4(p_6_in[9]),
        .I5(\r[irl][3][2]_i_18_n_0 ),
        .O(\r[irl][3][0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000F4FFFF00F4)) 
    \r[irl][3][0]_i_7 
       (.I0(\r[irl][3][2]_i_14_n_0 ),
        .I1(\r[irl][3][3]_i_11_n_0 ),
        .I2(\r[irl][3][3]_i_18_n_0 ),
        .I3(\r[irl][3][3]_i_19_n_0 ),
        .I4(\r[irl][3][2]_i_12_n_0 ),
        .I5(\r[irl][3][0]_i_9_n_0 ),
        .O(\r[irl][3][0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF000C00FF000E00)) 
    \r[irl][3][0]_i_8 
       (.I0(\r[irl][3][3]_i_13_n_0 ),
        .I1(\r[irl][3][2]_i_9_n_0 ),
        .I2(\r[irl][3][2]_i_8_n_0 ),
        .I3(\r[irl][3][2]_i_7_n_0 ),
        .I4(\r[irl][3][2]_i_6_n_0 ),
        .I5(\r[irl][3][3]_i_14_n_0 ),
        .O(\r[irl][3][0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF00A800A800A8)) 
    \r[irl][3][0]_i_9 
       (.I0(\r_reg[imask][3]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[iforce][3]__0 [14]),
        .I3(p_6_in[15]),
        .I4(\r[irl][3][3]_i_22_n_0 ),
        .I5(\r[irl][3][3]_i_20_n_0 ),
        .O(\r[irl][3][0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDDDD0000DDDD000F)) 
    \r[irl][3][1]_i_1 
       (.I0(\r[irl][3][2]_i_3_n_0 ),
        .I1(\r[irl][3][1]_i_2_n_0 ),
        .I2(\r[irl][3][1]_i_3_n_0 ),
        .I3(\r[irl][3][1]_i_4_n_0 ),
        .I4(\r[irl][3][1]_i_5_n_0 ),
        .I5(\r[irl][3][1]_i_6_n_0 ),
        .O(\r[irl][3][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF100)) 
    \r[irl][3][1]_i_10 
       (.I0(\r[irl][3][1]_i_14_n_0 ),
        .I1(p_6_in[11]),
        .I2(\r[irl][3][3]_i_18_n_0 ),
        .I3(\r[irl][3][1]_i_17_n_0 ),
        .I4(\r[irl][3][1]_i_18_n_0 ),
        .O(\r[irl][3][1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][1]_i_11 
       (.I0(\r_reg[imask][3]__0 [3]),
        .I1(p_5_in[4]),
        .I2(\r_reg[iforce][3]__0 [3]),
        .O(\r[irl][3][1]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0E000E000E000000)) 
    \r[irl][3][1]_i_12 
       (.I0(\r[irl][3][2]_i_18_n_0 ),
        .I1(p_6_in[9]),
        .I2(\r[irl][3][3]_i_12_n_0 ),
        .I3(\r[irl][3][2]_i_15_n_0 ),
        .I4(\r[irl][3][1]_i_19_n_0 ),
        .I5(p_6_in[6]),
        .O(\r[irl][3][1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][1]_i_13 
       (.I0(p_6_in[3]),
        .I1(\r_reg[iforce][3]__0 [2]),
        .I2(p_5_in[3]),
        .I3(\r_reg[imask][3]__0 [2]),
        .O(\r[irl][3][1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][1]_i_14 
       (.I0(\r_reg[imask][3]__0 [10]),
        .I1(p_5_in[11]),
        .I2(\r_reg[iforce][3]__0 [10]),
        .O(\r[irl][3][1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFA800)) 
    \r[irl][3][1]_i_15 
       (.I0(\r_reg[imask][3]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][3]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][3][2]_i_8_n_0 ),
        .O(\r[irl][3][1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000777F)) 
    \r[irl][3][1]_i_16 
       (.I0(p_6_in[15]),
        .I1(\r_reg[imask][3]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[iforce][3]__0 [14]),
        .I4(\r[irl][3][2]_i_6_n_0 ),
        .O(\r[irl][3][1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FF57)) 
    \r[irl][3][1]_i_17 
       (.I0(\r_reg[imask][3]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][3]__0 [11]),
        .I3(p_6_in[12]),
        .I4(\r[irl][3][3]_i_22_n_0 ),
        .O(\r[irl][3][1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00A8FFFF)) 
    \r[irl][3][1]_i_18 
       (.I0(\r_reg[imask][3]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[iforce][3]__0 [14]),
        .I3(p_6_in[15]),
        .I4(\r[irl][3][3]_i_20_n_0 ),
        .O(\r[irl][3][1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][1]_i_19 
       (.I0(\r_reg[imask][3]__0 [5]),
        .I1(p_5_in[6]),
        .I2(\r_reg[iforce][3]__0 [5]),
        .O(\r[irl][3][1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00F4F4)) 
    \r[irl][3][1]_i_2 
       (.I0(\r[irl][3][1]_i_7_n_0 ),
        .I1(p_6_in[7]),
        .I2(\r[irl][3][1]_i_8_n_0 ),
        .I3(\r[irl][3][1]_i_9_n_0 ),
        .I4(\r[irl][3][3]_i_2_n_0 ),
        .O(\r[irl][3][1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF2222000F2222)) 
    \r[irl][3][1]_i_3 
       (.I0(\r[irl][3][3]_i_4_n_0 ),
        .I1(\r[irl][3][1]_i_10_n_0 ),
        .I2(p_6_in[4]),
        .I3(\r[irl][3][1]_i_11_n_0 ),
        .I4(\r[irl][3][1]_i_12_n_0 ),
        .I5(\r[irl][3][2]_i_13_n_0 ),
        .O(\r[irl][3][1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][1]_i_4 
       (.I0(p_6_in[1]),
        .I1(\r_reg[iforce][3]__0 [0]),
        .I2(p_5_in[1]),
        .I3(\r_reg[imask][3]__0 [0]),
        .O(\r[irl][3][1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF2FF)) 
    \r[irl][3][1]_i_5 
       (.I0(p_6_in[3]),
        .I1(\r[irl][3][3]_i_10_n_0 ),
        .I2(\r[irl][3][3]_i_9_n_0 ),
        .I3(\r[irl][3][3]_i_8_n_0 ),
        .I4(\r[irl][3][3]_i_7_n_0 ),
        .O(\r[irl][3][1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FF570000)) 
    \r[irl][3][1]_i_6 
       (.I0(\r_reg[imask][3]__0 [1]),
        .I1(p_5_in[2]),
        .I2(\r_reg[iforce][3]__0 [1]),
        .I3(p_6_in[2]),
        .I4(\r[irl][3][2]_i_5_n_0 ),
        .I5(\r[irl][3][1]_i_13_n_0 ),
        .O(\r[irl][3][1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][1]_i_7 
       (.I0(\r_reg[imask][3]__0 [6]),
        .I1(p_5_in[7]),
        .I2(\r_reg[iforce][3]__0 [6]),
        .O(\r[irl][3][1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][1]_i_8 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][3]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][3]__0 [5]),
        .O(\r[irl][3][1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00F4FFFF)) 
    \r[irl][3][1]_i_9 
       (.I0(\r[irl][3][1]_i_14_n_0 ),
        .I1(p_6_in[11]),
        .I2(\r[irl][3][3]_i_13_n_0 ),
        .I3(\r[irl][3][1]_i_15_n_0 ),
        .I4(\r[irl][3][1]_i_16_n_0 ),
        .O(\r[irl][3][1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7070707070FF7070)) 
    \r[irl][3][2]_i_1 
       (.I0(\r[irl][3][2]_i_2_n_0 ),
        .I1(\r[irl][3][3]_i_2_n_0 ),
        .I2(\r[irl][3][2]_i_3_n_0 ),
        .I3(\r[irl][3][2]_i_4_n_0 ),
        .I4(\r[irl][3][3]_i_3_n_0 ),
        .I5(\r[irl][3][2]_i_5_n_0 ),
        .O(\r[irl][3][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFEFEFFFE)) 
    \r[irl][3][2]_i_10 
       (.I0(\r[irl][3][1]_i_8_n_0 ),
        .I1(\r[irl][3][3]_i_16_n_0 ),
        .I2(\r[irl][3][3]_i_5_n_0 ),
        .I3(p_6_in[9]),
        .I4(\r[irl][3][2]_i_18_n_0 ),
        .I5(\r[irl][3][3]_i_6_n_0 ),
        .O(\r[irl][3][2]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF00A8)) 
    \r[irl][3][2]_i_11 
       (.I0(\r_reg[imask][3]__0 [8]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][3]__0 [8]),
        .I3(p_6_in[9]),
        .I4(\r[irl][3][3]_i_12_n_0 ),
        .O(\r[irl][3][2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFDFDFDFF)) 
    \r[irl][3][2]_i_12 
       (.I0(\r[irl][3][3]_i_20_n_0 ),
        .I1(\r[irl][3][3]_i_21_n_0 ),
        .I2(\r[irl][3][3]_i_22_n_0 ),
        .I3(p_6_in[12]),
        .I4(\r[irl][3][2]_i_19_n_0 ),
        .O(\r[irl][3][2]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][2]_i_13 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][3]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][3]__0 [4]),
        .O(\r[irl][3][2]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][2]_i_14 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][3]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][3]__0 [8]),
        .O(\r[irl][3][2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55551115)) 
    \r[irl][3][2]_i_15 
       (.I0(\r[irl][3][3]_i_11_n_0 ),
        .I1(\r_reg[imask][3]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[iforce][3]__0 [6]),
        .I4(p_6_in[7]),
        .O(\r[irl][3][2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][2]_i_16 
       (.I0(p_6_in[6]),
        .I1(\r_reg[iforce][3]__0 [5]),
        .I2(p_5_in[6]),
        .I3(\r_reg[imask][3]__0 [5]),
        .O(\r[irl][3][2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][2]_i_17 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][3]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][3]__0 [3]),
        .O(\r[irl][3][2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][2]_i_18 
       (.I0(\r_reg[imask][3]__0 [8]),
        .I1(p_5_in[9]),
        .I2(\r_reg[iforce][3]__0 [8]),
        .O(\r[irl][3][2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][2]_i_19 
       (.I0(\r_reg[imask][3]__0 [11]),
        .I1(p_5_in[12]),
        .I2(\r_reg[iforce][3]__0 [11]),
        .O(\r[irl][3][2]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \r[irl][3][2]_i_2 
       (.I0(\r[irl][3][2]_i_6_n_0 ),
        .I1(\r[irl][3][2]_i_7_n_0 ),
        .I2(\r[irl][3][2]_i_8_n_0 ),
        .I3(\r[irl][3][2]_i_9_n_0 ),
        .O(\r[irl][3][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][3][2]_i_3 
       (.I0(\r[irl][3][3]_i_9_n_0 ),
        .I1(p_6_in[5]),
        .I2(\r_reg[iforce][3]__0 [4]),
        .I3(p_5_in[5]),
        .I4(\r_reg[imask][3]__0 [4]),
        .I5(\r[irl][3][2]_i_10_n_0 ),
        .O(\r[irl][3][2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000BBBAAAAA)) 
    \r[irl][3][2]_i_4 
       (.I0(\r[irl][3][2]_i_11_n_0 ),
        .I1(p_6_in[8]),
        .I2(\r_reg[iforce][3]__0 [7]),
        .I3(p_5_in[8]),
        .I4(\r_reg[imask][3]__0 [7]),
        .I5(\r[irl][3][2]_i_12_n_0 ),
        .O(\r[irl][3][2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \r[irl][3][2]_i_5 
       (.I0(\r[irl][3][2]_i_13_n_0 ),
        .I1(\r[irl][3][2]_i_14_n_0 ),
        .I2(\r[irl][3][3]_i_12_n_0 ),
        .I3(\r[irl][3][2]_i_15_n_0 ),
        .I4(\r[irl][3][2]_i_16_n_0 ),
        .I5(\r[irl][3][2]_i_17_n_0 ),
        .O(\r[irl][3][2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][2]_i_6 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][3]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][3]__0 [13]),
        .O(\r[irl][3][2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1FFF)) 
    \r[irl][3][2]_i_7 
       (.I0(\r_reg[iforce][3]__0 [14]),
        .I1(p_5_in[15]),
        .I2(\r_reg[imask][3]__0 [14]),
        .I3(p_6_in[15]),
        .O(\r[irl][3][2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][2]_i_8 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][3]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][3]__0 [12]),
        .O(\r[irl][3][2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][2]_i_9 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][3]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][3]__0 [11]),
        .O(\r[irl][3][2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \r[irl][3][3]_i_1 
       (.I0(\r[irl][3][3]_i_2_n_0 ),
        .I1(\r[irl][3][3]_i_3_n_0 ),
        .I2(\r[irl][3][3]_i_4_n_0 ),
        .O(\r[irl][3][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h57)) 
    \r[irl][3][3]_i_10 
       (.I0(\r_reg[imask][3]__0 [2]),
        .I1(p_5_in[3]),
        .I2(\r_reg[iforce][3]__0 [2]),
        .O(\r[irl][3][3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_11 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][3]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][3]__0 [7]),
        .O(\r[irl][3][3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFEF)) 
    \r[irl][3][3]_i_12 
       (.I0(\r[irl][3][3]_i_18_n_0 ),
        .I1(\r[irl][3][3]_i_19_n_0 ),
        .I2(\r[irl][3][3]_i_20_n_0 ),
        .I3(\r[irl][3][3]_i_21_n_0 ),
        .I4(\r[irl][3][3]_i_22_n_0 ),
        .I5(\r[irl][3][3]_i_23_n_0 ),
        .O(\r[irl][3][3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_13 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][3]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][3]__0 [9]),
        .O(\r[irl][3][3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_14 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][3]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][3]__0 [10]),
        .O(\r[irl][3][3]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_15 
       (.I0(p_6_in[9]),
        .I1(\r_reg[iforce][3]__0 [8]),
        .I2(p_5_in[9]),
        .I3(\r_reg[imask][3]__0 [8]),
        .O(\r[irl][3][3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_16 
       (.I0(p_6_in[7]),
        .I1(\r_reg[iforce][3]__0 [6]),
        .I2(p_5_in[7]),
        .I3(\r_reg[imask][3]__0 [6]),
        .O(\r[irl][3][3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_17 
       (.I0(p_6_in[5]),
        .I1(\r_reg[iforce][3]__0 [4]),
        .I2(p_5_in[5]),
        .I3(\r_reg[imask][3]__0 [4]),
        .O(\r[irl][3][3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_18 
       (.I0(p_6_in[10]),
        .I1(\r_reg[iforce][3]__0 [9]),
        .I2(p_5_in[10]),
        .I3(\r_reg[imask][3]__0 [9]),
        .O(\r[irl][3][3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_19 
       (.I0(p_6_in[11]),
        .I1(\r_reg[iforce][3]__0 [10]),
        .I2(p_5_in[11]),
        .I3(\r_reg[imask][3]__0 [10]),
        .O(\r[irl][3][3]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFEEEAAAAA)) 
    \r[irl][3][3]_i_2 
       (.I0(\r[irl][3][3]_i_5_n_0 ),
        .I1(p_6_in[9]),
        .I2(\r_reg[iforce][3]__0 [8]),
        .I3(p_5_in[9]),
        .I4(\r_reg[imask][3]__0 [8]),
        .I5(\r[irl][3][3]_i_6_n_0 ),
        .O(\r[irl][3][3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hABFF)) 
    \r[irl][3][3]_i_20 
       (.I0(p_6_in[14]),
        .I1(\r_reg[iforce][3]__0 [13]),
        .I2(p_5_in[14]),
        .I3(\r_reg[imask][3]__0 [13]),
        .O(\r[irl][3][3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_21 
       (.I0(p_6_in[15]),
        .I1(\r_reg[iforce][3]__0 [14]),
        .I2(p_5_in[15]),
        .I3(\r_reg[imask][3]__0 [14]),
        .O(\r[irl][3][3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_22 
       (.I0(p_6_in[13]),
        .I1(\r_reg[iforce][3]__0 [12]),
        .I2(p_5_in[13]),
        .I3(\r_reg[imask][3]__0 [12]),
        .O(\r[irl][3][3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5400)) 
    \r[irl][3][3]_i_23 
       (.I0(p_6_in[12]),
        .I1(\r_reg[iforce][3]__0 [11]),
        .I2(p_5_in[12]),
        .I3(\r_reg[imask][3]__0 [11]),
        .O(\r[irl][3][3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000004000404)) 
    \r[irl][3][3]_i_3 
       (.I0(\r[irl][3][3]_i_7_n_0 ),
        .I1(\r[irl][3][3]_i_8_n_0 ),
        .I2(\r[irl][3][3]_i_9_n_0 ),
        .I3(\r[irl][3][3]_i_10_n_0 ),
        .I4(p_6_in[3]),
        .I5(\r[irl][3][1]_i_4_n_0 ),
        .O(\r[irl][3][3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEFEFEEEEEEEEEE)) 
    \r[irl][3][3]_i_4 
       (.I0(\r[irl][3][3]_i_11_n_0 ),
        .I1(\r[irl][3][3]_i_12_n_0 ),
        .I2(p_6_in[9]),
        .I3(\r_reg[iforce][3]__0 [8]),
        .I4(p_5_in[9]),
        .I5(\r_reg[imask][3]__0 [8]),
        .O(\r[irl][3][3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_5 
       (.I0(p_6_in[8]),
        .I1(\r_reg[iforce][3]__0 [7]),
        .I2(p_5_in[8]),
        .I3(\r_reg[imask][3]__0 [7]),
        .O(\r[irl][3][3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFEFF)) 
    \r[irl][3][3]_i_6 
       (.I0(\r[irl][3][3]_i_13_n_0 ),
        .I1(\r[irl][3][3]_i_14_n_0 ),
        .I2(\r[irl][3][2]_i_6_n_0 ),
        .I3(\r[irl][3][2]_i_7_n_0 ),
        .I4(\r[irl][3][2]_i_8_n_0 ),
        .I5(\r[irl][3][2]_i_9_n_0 ),
        .O(\r[irl][3][3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_7 
       (.I0(p_6_in[2]),
        .I1(\r_reg[iforce][3]__0 [1]),
        .I2(p_5_in[2]),
        .I3(\r_reg[imask][3]__0 [1]),
        .O(\r[irl][3][3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \r[irl][3][3]_i_8 
       (.I0(\r[irl][3][3]_i_6_n_0 ),
        .I1(\r[irl][3][3]_i_15_n_0 ),
        .I2(\r[irl][3][3]_i_5_n_0 ),
        .I3(\r[irl][3][3]_i_16_n_0 ),
        .I4(\r[irl][3][1]_i_8_n_0 ),
        .I5(\r[irl][3][3]_i_17_n_0 ),
        .O(\r[irl][3][3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA800)) 
    \r[irl][3][3]_i_9 
       (.I0(p_6_in[4]),
        .I1(\r_reg[iforce][3]__0 [3]),
        .I2(p_5_in[4]),
        .I3(\r_reg[imask][3]__0 [3]),
        .O(\r[irl][3][3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4444444444444445)) 
    \r[newaddr][2]_i_1 
       (.I0(v),
        .I1(\irqo[3][pwdnewaddr] [2]),
        .I2(r_reg),
        .I3(\r_reg[clkcount_n_0_][1] ),
        .I4(\r_reg[clkcount_n_0_][2] ),
        .I5(\r[newaddr][2]_i_2_n_0 ),
        .O(\r[newaddr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \r[newaddr][2]_i_2 
       (.I0(\irqo[1][svtclrtt] ),
        .I1(\irqo[0][svtclrtt] ),
        .I2(\irqo[2][svtclrtt] ),
        .I3(\irqo[3][svtclrtt] ),
        .O(\r[newaddr][2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800000000000)) 
    \r[newaddr][31]_i_1 
       (.I0(\apbi[pwrite] ),
        .I1(\apbi[penable] ),
        .I2(apbi[2]),
        .I3(\apbi[paddr] [5]),
        .I4(\apbi[paddr] [7]),
        .I5(\apbi[paddr] [6]),
        .O(v));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r[setaddr][0]_i_1 
       (.I0(rst),
        .O(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555D0000000C)) 
    \r[setaddr][0]_i_2 
       (.I0(\r[setaddr][0]_i_3_n_0 ),
        .I1(v),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\irqo[0][svtclrtt] ),
        .O(\r[setaddr][0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000FFFE0000)) 
    \r[setaddr][0]_i_3 
       (.I0(\irqo[3][svtclrtt] ),
        .I1(\irqo[2][svtclrtt] ),
        .I2(\irqo[0][svtclrtt] ),
        .I3(\irqo[1][svtclrtt] ),
        .I4(\irqo[3][pwdnewaddr] [2]),
        .I5(\r[forceerr][0]_i_2_n_0 ),
        .O(\r[setaddr][0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h55555D5500000C00)) 
    \r[setaddr][1]_i_1 
       (.I0(\r[setaddr][0]_i_3_n_0 ),
        .I1(v),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\irqo[1][svtclrtt] ),
        .O(\r[setaddr][1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5575555500300000)) 
    \r[setaddr][2]_i_1 
       (.I0(\r[setaddr][0]_i_3_n_0 ),
        .I1(\apbi[paddr] [2]),
        .I2(\apbi[paddr] [3]),
        .I3(\apbi[paddr] [4]),
        .I4(v),
        .I5(\irqo[2][svtclrtt] ),
        .O(\r[setaddr][2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5D5555550C000000)) 
    \r[setaddr][3]_i_1 
       (.I0(\r[setaddr][0]_i_3_n_0 ),
        .I1(v),
        .I2(\apbi[paddr] [4]),
        .I3(\apbi[paddr] [2]),
        .I4(\apbi[paddr] [3]),
        .I5(\irqo[3][svtclrtt] ),
        .O(\r[setaddr][3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFB08)) 
    \r[setaddrboot]_i_1 
       (.I0(\apbi[pwdata] [0]),
        .I1(v),
        .I2(\apbi[paddr] [4]),
        .I3(\r_reg[setaddrboot_n_0_] ),
        .O(\r[setaddrboot]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[clkcount][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(r),
        .Q(r_reg),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[clkcount][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[clkcount][1]_i_1_n_0 ),
        .Q(\r_reg[clkcount_n_0_][1] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[clkcount][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[clkcount][2]_i_1_n_0 ),
        .Q(\r_reg[clkcount_n_0_][2] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[cpurst][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\v[cpurst]1_out [0]),
        .Q(\irqo[0][resume] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[cpurst][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\v[cpurst]1_out [1]),
        .Q(\irqo[1][resume] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[cpurst][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\v[cpurst]1_out [2]),
        .Q(\irqo[2][resume] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[cpurst][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\v[cpurst]1_out [3]),
        .Q(\irqo[3][resume] ),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[forceerr][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[forceerr][0]_i_1_n_0 ),
        .Q(\irqo[0][forceerr] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[forceerr][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[forceerr][1]_i_1_n_0 ),
        .Q(\irqo[1][forceerr] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[forceerr][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[forceerr][2]_i_1_n_0 ),
        .Q(\irqo[2][forceerr] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[forceerr][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[forceerr][3]_i_1_n_0 ),
        .Q(\irqo[3][forceerr] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][10] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [10]),
        .Q(p_0_in14_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][11] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [11]),
        .Q(p_0_in12_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][12] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [12]),
        .Q(p_0_in10_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][13] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [13]),
        .Q(p_0_in8_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][14] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [14]),
        .Q(p_0_in6_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][15] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [15]),
        .Q(p_0_in4_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][1] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [1]),
        .Q(\r_reg[ibroadcast_n_0_][1] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][2] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [2]),
        .Q(p_0_in30_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][3] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [3]),
        .Q(p_0_in28_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][4] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [4]),
        .Q(p_0_in26_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][5] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [5]),
        .Q(p_0_in24_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][6] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [6]),
        .Q(p_0_in22_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][7] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [7]),
        .Q(p_0_in20_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][8] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [8]),
        .Q(p_0_in18_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ibroadcast][9] 
       (.C(clk),
        .CE(\v[ibroadcast] ),
        .D(\apbi[pwdata] [9]),
        .Q(p_0_in16_in),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][10] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][10]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][11] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][11]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][12] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][12]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][13] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][13]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][14] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][14]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][15] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][15]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][1]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][2]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][3]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][4] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][4]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][5] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][5]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][6] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][6]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][7] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][7]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][8] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][8]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][0][9] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][0][9]_i_1_n_0 ),
        .Q(\r_reg[iforce][0]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][10] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][10]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][11] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][11]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][12] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][12]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][13] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][13]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][14] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][14]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][15] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][15]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][1]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][2]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][3]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][4] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][4]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][5] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][5]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][6] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][6]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][7] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][7]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][8] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][8]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][1][9] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][1][9]_i_1_n_0 ),
        .Q(\r_reg[iforce][1]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][10] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][10]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][11] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][11]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][12] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][12]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][13] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][13]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][14] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][14]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][15] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][15]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][1]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][2]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][3]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][4] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][4]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][5] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][5]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][6] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][6]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][7] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][7]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][8] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][8]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][2][9] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][2][9]_i_1_n_0 ),
        .Q(\r_reg[iforce][2]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][10] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][10]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][11] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][11]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][12] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][12]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][13] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][13]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][14] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][14]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][15] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][15]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][1]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][2]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][3]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][4] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][4]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][5] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][5]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][6] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][6]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][7] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][7]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][8] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][8]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[iforce][3][9] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[iforce][3][9]_i_1_n_0 ),
        .Q(\r_reg[iforce][3]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][10] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [10]),
        .Q(p_6_in[10]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][11] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [11]),
        .Q(p_6_in[11]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][12] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [12]),
        .Q(p_6_in[12]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][13] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [13]),
        .Q(p_6_in[13]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][14] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [14]),
        .Q(p_6_in[14]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][15] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [15]),
        .Q(p_6_in[15]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][1] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [1]),
        .Q(p_6_in[1]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][2] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [2]),
        .Q(p_6_in[2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][3] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [3]),
        .Q(p_6_in[3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][4] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [4]),
        .Q(p_6_in[4]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][5] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [5]),
        .Q(p_6_in[5]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][6] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [6]),
        .Q(p_6_in[6]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][7] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [7]),
        .Q(p_6_in[7]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][8] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [8]),
        .Q(p_6_in[8]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ilevel][9] 
       (.C(clk),
        .CE(\v[ilevel] ),
        .D(\apbi[pwdata] [9]),
        .Q(p_6_in[9]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][10] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [10]),
        .Q(\r_reg[imask][0]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][11] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [11]),
        .Q(\r_reg[imask][0]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][12] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [12]),
        .Q(\r_reg[imask][0]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][13] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [13]),
        .Q(\r_reg[imask][0]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][14] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [14]),
        .Q(\r_reg[imask][0]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][15] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [15]),
        .Q(\r_reg[imask][0]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][1] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [1]),
        .Q(\r_reg[imask][0]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][2] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [2]),
        .Q(\r_reg[imask][0]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][3] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [3]),
        .Q(\r_reg[imask][0]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][4] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [4]),
        .Q(\r_reg[imask][0]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][5] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [5]),
        .Q(\r_reg[imask][0]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][6] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [6]),
        .Q(\r_reg[imask][0]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][7] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [7]),
        .Q(\r_reg[imask][0]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][8] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [8]),
        .Q(\r_reg[imask][0]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][0][9] 
       (.C(clk),
        .CE(\v[imask][0] ),
        .D(\apbi[pwdata] [9]),
        .Q(\r_reg[imask][0]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][10] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [10]),
        .Q(\r_reg[imask][1]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][11] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [11]),
        .Q(\r_reg[imask][1]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][12] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [12]),
        .Q(\r_reg[imask][1]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][13] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [13]),
        .Q(\r_reg[imask][1]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][14] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [14]),
        .Q(\r_reg[imask][1]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][15] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [15]),
        .Q(\r_reg[imask][1]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][1] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [1]),
        .Q(\r_reg[imask][1]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][2] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [2]),
        .Q(\r_reg[imask][1]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][3] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [3]),
        .Q(\r_reg[imask][1]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][4] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [4]),
        .Q(\r_reg[imask][1]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][5] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [5]),
        .Q(\r_reg[imask][1]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][6] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [6]),
        .Q(\r_reg[imask][1]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][7] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [7]),
        .Q(\r_reg[imask][1]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][8] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [8]),
        .Q(\r_reg[imask][1]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][1][9] 
       (.C(clk),
        .CE(\v[imask][1] ),
        .D(\apbi[pwdata] [9]),
        .Q(\r_reg[imask][1]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][10] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [10]),
        .Q(\r_reg[imask][2]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][11] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [11]),
        .Q(\r_reg[imask][2]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][12] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [12]),
        .Q(\r_reg[imask][2]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][13] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [13]),
        .Q(\r_reg[imask][2]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][14] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [14]),
        .Q(\r_reg[imask][2]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][15] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [15]),
        .Q(\r_reg[imask][2]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][1] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [1]),
        .Q(\r_reg[imask][2]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][2] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [2]),
        .Q(\r_reg[imask][2]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][3] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [3]),
        .Q(\r_reg[imask][2]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][4] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [4]),
        .Q(\r_reg[imask][2]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][5] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [5]),
        .Q(\r_reg[imask][2]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][6] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [6]),
        .Q(\r_reg[imask][2]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][7] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [7]),
        .Q(\r_reg[imask][2]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][8] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [8]),
        .Q(\r_reg[imask][2]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][2][9] 
       (.C(clk),
        .CE(\v[imask][2] ),
        .D(\apbi[pwdata] [9]),
        .Q(\r_reg[imask][2]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][10] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [10]),
        .Q(\r_reg[imask][3]__0 [9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][11] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [11]),
        .Q(\r_reg[imask][3]__0 [10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][12] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [12]),
        .Q(\r_reg[imask][3]__0 [11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][13] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [13]),
        .Q(\r_reg[imask][3]__0 [12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][14] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [14]),
        .Q(\r_reg[imask][3]__0 [13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][15] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [15]),
        .Q(\r_reg[imask][3]__0 [14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][1] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [1]),
        .Q(\r_reg[imask][3]__0 [0]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][2] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [2]),
        .Q(\r_reg[imask][3]__0 [1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][3] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [3]),
        .Q(\r_reg[imask][3]__0 [2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][4] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [4]),
        .Q(\r_reg[imask][3]__0 [3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][5] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [5]),
        .Q(\r_reg[imask][3]__0 [4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][6] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [6]),
        .Q(\r_reg[imask][3]__0 [5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][7] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [7]),
        .Q(\r_reg[imask][3]__0 [6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][8] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [8]),
        .Q(\r_reg[imask][3]__0 [7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[imask][3][9] 
       (.C(clk),
        .CE(\v[imask][3] ),
        .D(\apbi[pwdata] [9]),
        .Q(\r_reg[imask][3]__0 [8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][10] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][10]_i_1_n_0 ),
        .Q(p_5_in[10]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][11] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][11]_i_1_n_0 ),
        .Q(p_5_in[11]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][12] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][12]_i_1_n_0 ),
        .Q(p_5_in[12]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][13] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][13]_i_1_n_0 ),
        .Q(p_5_in[13]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][14] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][14]_i_1_n_0 ),
        .Q(p_5_in[14]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][15] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][15]_i_1_n_0 ),
        .Q(p_5_in[15]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][1]_i_1_n_0 ),
        .Q(p_5_in[1]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][2]_i_1_n_0 ),
        .Q(p_5_in[2]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][3]_i_1_n_0 ),
        .Q(p_5_in[3]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][4] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][4]_i_1_n_0 ),
        .Q(p_5_in[4]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][5] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][5]_i_1_n_0 ),
        .Q(p_5_in[5]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][6] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][6]_i_1_n_0 ),
        .Q(p_5_in[6]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][7] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][7]_i_1_n_0 ),
        .Q(p_5_in[7]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][8] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][8]_i_1_n_0 ),
        .Q(p_5_in[8]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[ipend][9] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[ipend][9]_i_1_n_0 ),
        .Q(p_5_in[9]),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][0][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][0][0]_i_1_n_0 ),
        .Q(\irqo[0][irl] [0]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][0][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][0][1]_i_1_n_0 ),
        .Q(\irqo[0][irl] [1]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][0][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][0][2]_i_1_n_0 ),
        .Q(\irqo[0][irl] [2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][0][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][0][3]_i_1_n_0 ),
        .Q(\irqo[0][irl] [3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][1][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][1][0]_i_1_n_0 ),
        .Q(\irqo[1][irl] [0]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][1][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][1][1]_i_1_n_0 ),
        .Q(\irqo[1][irl] [1]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][1][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][1][2]_i_1_n_0 ),
        .Q(\irqo[1][irl] [2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][1][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][1][3]_i_1_n_0 ),
        .Q(\irqo[1][irl] [3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][2][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][2][0]_i_1_n_0 ),
        .Q(\irqo[2][irl] [0]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][2][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][2][1]_i_1_n_0 ),
        .Q(\irqo[2][irl] [1]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][2][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][2][2]_i_1_n_0 ),
        .Q(\irqo[2][irl] [2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][2][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][2][3]_i_1_n_0 ),
        .Q(\irqo[2][irl] [3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][3][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][3][0]_i_1_n_0 ),
        .Q(\irqo[3][irl] [0]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][3][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][3][1]_i_1_n_0 ),
        .Q(\irqo[3][irl] [1]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][3][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][3][2]_i_1_n_0 ),
        .Q(\irqo[3][irl] [2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[irl][3][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[irl][3][3]_i_1_n_0 ),
        .Q(\irqo[3][irl] [3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][10] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [10]),
        .Q(\irqo[3][pwdnewaddr] [10]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][11] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [11]),
        .Q(\irqo[3][pwdnewaddr] [11]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][12] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [12]),
        .Q(\irqo[3][pwdnewaddr] [12]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][13] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [13]),
        .Q(\irqo[3][pwdnewaddr] [13]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][14] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [14]),
        .Q(\irqo[3][pwdnewaddr] [14]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][15] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [15]),
        .Q(\irqo[3][pwdnewaddr] [15]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][16] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [16]),
        .Q(\irqo[3][pwdnewaddr] [16]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][17] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [17]),
        .Q(\irqo[3][pwdnewaddr] [17]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][18] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [18]),
        .Q(\irqo[3][pwdnewaddr] [18]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][19] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [19]),
        .Q(\irqo[3][pwdnewaddr] [19]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][20] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [20]),
        .Q(\irqo[3][pwdnewaddr] [20]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][21] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [21]),
        .Q(\irqo[3][pwdnewaddr] [21]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][22] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [22]),
        .Q(\irqo[3][pwdnewaddr] [22]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][23] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [23]),
        .Q(\irqo[3][pwdnewaddr] [23]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][24] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [24]),
        .Q(\irqo[3][pwdnewaddr] [24]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][25] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [25]),
        .Q(\irqo[3][pwdnewaddr] [25]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][26] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [26]),
        .Q(\irqo[3][pwdnewaddr] [26]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][27] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [27]),
        .Q(\irqo[3][pwdnewaddr] [27]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][28] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [28]),
        .Q(\irqo[3][pwdnewaddr] [28]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][29] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [29]),
        .Q(\irqo[3][pwdnewaddr] [29]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[newaddr][2]_i_1_n_0 ),
        .Q(\irqo[3][pwdnewaddr] [2]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][30] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [30]),
        .Q(\irqo[3][pwdnewaddr] [30]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][31] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [31]),
        .Q(\irqo[3][pwdnewaddr] [31]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][3] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [3]),
        .Q(\irqo[3][pwdnewaddr] [3]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][4] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [4]),
        .Q(\irqo[3][pwdnewaddr] [4]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][5] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [5]),
        .Q(\irqo[3][pwdnewaddr] [5]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][6] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [6]),
        .Q(\irqo[3][pwdnewaddr] [6]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][7] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [7]),
        .Q(\irqo[3][pwdnewaddr] [7]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][8] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [8]),
        .Q(\irqo[3][pwdnewaddr] [8]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[newaddr][9] 
       (.C(clk),
        .CE(v),
        .D(\apbi[pwdata] [9]),
        .Q(\irqo[3][pwdnewaddr] [9]),
        .R(irqo));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[setaddr][0] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[setaddr][0]_i_2_n_0 ),
        .Q(\irqo[0][svtclrtt] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[setaddr][1] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[setaddr][1]_i_1_n_0 ),
        .Q(\irqo[1][svtclrtt] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[setaddr][2] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[setaddr][2]_i_1_n_0 ),
        .Q(\irqo[2][svtclrtt] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[setaddr][3] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[setaddr][3]_i_1_n_0 ),
        .Q(\irqo[3][svtclrtt] ),
        .R(p_0_in));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_reg[setaddrboot] 
       (.C(clk),
        .CE(\^irqo[3][index] ),
        .D(\r[setaddrboot]_i_1_n_0 ),
        .Q(\r_reg[setaddrboot_n_0_] ),
        .R(irqo));
endmodule
