module sha3_low_throughput
   (clk,
    reset,
    in,
    in_ready,
    is_last,
    byte_num,
    buffer_full,
    out,
    backdoor,
    out_ready);
  output backdoor;
  input clk;
  input reset;
  input [31:0]in;
  input in_ready;
  input is_last;
  input [1:0]byte_num;
  output buffer_full;
  output [511:0]out;
  output out_ready;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire buffer_full;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1:0]byte_num;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire done_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/calc ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/calc0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/i_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1000] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1001] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1002] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1003] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1004] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1005] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1006] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1007] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1008] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1009] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[100] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1010] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1011] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1012] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1013] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1014] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1015] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1016] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1017] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1018] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1019] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[101] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1020] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1021] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1022] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1023] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1024] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1025] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1026] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1027] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1028] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1029] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[102] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1030] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1031] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1032] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1033] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1034] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1035] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1036] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1037] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1038] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1039] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[103] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1040] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1041] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1042] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1043] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1044] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1045] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1046] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1047] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1048] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1049] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[104] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1050] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1051] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1052] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1053] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1054] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1055] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1056] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1057] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1058] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1059] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[105] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1060] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1061] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1062] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1063] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1064] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1065] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1066] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1067] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1068] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1069] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[106] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1070] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1071] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1072] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1073] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1074] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1075] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1076] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1077] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1078] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1079] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[107] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1080] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1081] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1082] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1083] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1084] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1085] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1086] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1087] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[108] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[109] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[110] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[111] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[112] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[113] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[114] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[115] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[116] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[117] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[118] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[119] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[120] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[121] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[122] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[123] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[124] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[125] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[126] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[127] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[128] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[129] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[130] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[131] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[132] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[133] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[134] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[135] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[136] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[137] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[138] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[139] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[140] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[141] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[142] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[143] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[144] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[145] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[146] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[147] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[148] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[149] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[150] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[151] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[152] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[153] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[154] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[155] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[156] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[157] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[158] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[159] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[160] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[161] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[162] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[163] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[164] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[165] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[166] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[167] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[168] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[169] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[170] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[171] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[172] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[173] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[174] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[175] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[176] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[177] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[178] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[179] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[180] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[181] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[182] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[183] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[184] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[185] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[186] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[187] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[188] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[189] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[190] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[191] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[192] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[193] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[194] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[195] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[196] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[197] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[198] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[199] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[200] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[201] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[202] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[203] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[204] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[205] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[206] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[207] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[208] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[209] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[210] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[211] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[212] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[213] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[214] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[215] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[216] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[217] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[218] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[219] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[220] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[221] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[222] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[223] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[224] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[225] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[226] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[227] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[228] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[229] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[230] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[231] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[232] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[233] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[234] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[235] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[236] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[237] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[238] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[239] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[240] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[241] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[242] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[243] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[244] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[245] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[246] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[247] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[248] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[249] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[250] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[251] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[252] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[253] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[254] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[255] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[256] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[257] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[258] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[259] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[260] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[261] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[262] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[263] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[264] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[265] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[266] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[267] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[268] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[269] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[270] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[271] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[272] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[273] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[274] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[275] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[276] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[277] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[278] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[279] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[280] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[281] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[282] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[283] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[284] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[285] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[286] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[287] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[288] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[289] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[290] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[291] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[292] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[293] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[294] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[295] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[296] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[297] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[298] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[299] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[300] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[301] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[302] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[303] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[304] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[305] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[306] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[307] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[308] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[309] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[310] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[311] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[312] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[313] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[314] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[315] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[316] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[317] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[318] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[319] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[320] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[321] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[322] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[323] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[324] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[325] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[326] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[327] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[328] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[329] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[330] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[331] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[332] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[333] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[334] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[335] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[336] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[337] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[338] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[339] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[340] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[341] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[342] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[343] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[344] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[345] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[346] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[347] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[348] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[349] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[350] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[351] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[352] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[353] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[354] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[355] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[356] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[357] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[358] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[359] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[360] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[361] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[362] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[363] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[364] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[365] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[366] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[367] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[368] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[369] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[370] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[371] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[372] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[373] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[374] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[375] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[376] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[377] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[378] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[379] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[380] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[381] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[382] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[383] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[384] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[385] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[386] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[387] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[388] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[389] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[390] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[391] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[392] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[393] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[394] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[395] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[396] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[397] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[398] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[399] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[400] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[401] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[402] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[403] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[404] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[405] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[406] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[407] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[408] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[409] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[410] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[411] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[412] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[413] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[414] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[415] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[416] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[417] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[418] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[419] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[420] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[421] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[422] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[423] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[424] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[425] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[426] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[427] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[428] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[429] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[430] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[431] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[432] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[433] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[434] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[435] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[436] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[437] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[438] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[439] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[440] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[441] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[442] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[443] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[444] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[445] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[446] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[447] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[448] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[449] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[450] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[451] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[452] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[453] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[454] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[455] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[456] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[457] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[458] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[459] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[460] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[461] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[462] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[463] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[464] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[465] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[466] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[467] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[468] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[469] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[470] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[471] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[472] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[473] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[474] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[475] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[476] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[477] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[478] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[479] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[480] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[481] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[482] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[483] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[484] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[485] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[486] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[487] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[488] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[489] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[490] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[491] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[492] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[493] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[494] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[495] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[496] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[497] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[498] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[499] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[500] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[501] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[502] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[503] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[504] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[505] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[506] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[507] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[508] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[509] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[510] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[511] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[512] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[513] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[514] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[515] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[516] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[517] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[518] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[519] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[520] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[521] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[522] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[523] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[524] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[525] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[526] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[527] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[528] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[529] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[530] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[531] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[532] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[533] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[534] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[535] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[536] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[537] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[538] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[539] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[540] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[541] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[542] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[543] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[544] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[545] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[546] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[547] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[548] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[549] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[550] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[551] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[552] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[553] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[554] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[555] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[556] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[557] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[558] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[559] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[560] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[561] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[562] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[563] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[564] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[565] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[566] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[567] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[568] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[569] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[570] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[571] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[572] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[573] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[574] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[575] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[576] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[577] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[578] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[579] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[580] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[581] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[582] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[583] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[584] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[585] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[586] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[587] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[588] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[589] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[590] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[591] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[592] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[593] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[594] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[595] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[596] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[597] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[598] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[599] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[600] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[601] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[602] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[603] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[604] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[605] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[606] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[607] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[608] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[609] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[610] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[611] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[612] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[613] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[614] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[615] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[616] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[617] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[618] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[619] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[620] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[621] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[622] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[623] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[624] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[625] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[626] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[627] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[628] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[629] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[630] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[631] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[632] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[633] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[634] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[635] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[636] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[637] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[638] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[639] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[640] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[641] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[642] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[643] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[644] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[645] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[646] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[647] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[648] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[649] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[64] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[650] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[651] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[652] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[653] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[654] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[655] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[656] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[657] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[658] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[659] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[65] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[660] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[661] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[662] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[663] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[664] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[665] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[666] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[667] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[668] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[669] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[66] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[670] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[671] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[672] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[673] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[674] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[675] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[676] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[677] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[678] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[679] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[67] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[680] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[681] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[682] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[683] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[684] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[685] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[686] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[687] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[688] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[689] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[68] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[690] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[691] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[692] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[693] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[694] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[695] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[696] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[697] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[698] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[699] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[69] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[700] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[701] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[702] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[703] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[704] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[705] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[706] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[707] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[708] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[709] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[70] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[710] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[711] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[712] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[713] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[714] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[715] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[716] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[717] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[718] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[719] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[71] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[720] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[721] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[722] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[723] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[724] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[725] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[726] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[727] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[728] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[729] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[72] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[730] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[731] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[732] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[733] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[734] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[735] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[736] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[737] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[738] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[739] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[73] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[740] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[741] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[742] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[743] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[744] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[745] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[746] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[747] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[748] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[749] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[74] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[750] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[751] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[752] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[753] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[754] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[755] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[756] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[757] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[758] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[759] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[75] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[760] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[761] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[762] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[763] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[764] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[765] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[766] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[767] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[768] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[769] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[76] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[770] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[771] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[772] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[773] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[774] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[775] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[776] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[777] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[778] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[779] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[77] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[780] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[781] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[782] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[783] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[784] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[785] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[786] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[787] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[788] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[789] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[78] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[790] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[791] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[792] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[793] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[794] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[795] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[796] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[797] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[798] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[799] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[79] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[800] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[801] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[802] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[803] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[804] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[805] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[806] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[807] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[808] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[809] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[80] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[810] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[811] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[812] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[813] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[814] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[815] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[816] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[817] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[818] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[819] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[81] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[820] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[821] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[822] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[823] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[824] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[825] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[826] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[827] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[828] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[829] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[82] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[830] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[831] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[832] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[833] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[834] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[835] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[836] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[837] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[838] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[839] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[83] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[840] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[841] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[842] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[843] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[844] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[845] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[846] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[847] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[848] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[849] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[84] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[850] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[851] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[852] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[853] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[854] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[855] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[856] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[857] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[858] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[859] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[85] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[860] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[861] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[862] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[863] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[864] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[865] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[866] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[867] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[868] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[869] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[86] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[870] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[871] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[872] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[873] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[874] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[875] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[876] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[877] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[878] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[879] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[87] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[880] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[881] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[882] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[883] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[884] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[885] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[886] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[887] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[888] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[889] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[88] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[890] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[891] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[892] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[893] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[894] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[895] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[896] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[897] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[898] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[899] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[89] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[900] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[901] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[902] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[903] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[904] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[905] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[906] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[907] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[908] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[909] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[90] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[910] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[911] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[912] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[913] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[914] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[915] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[916] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[917] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[918] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[919] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[91] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[920] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[921] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[922] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[923] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[924] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[925] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[926] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[927] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[928] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[929] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[92] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[930] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[931] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[932] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[933] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[934] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[935] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[936] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[937] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[938] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[939] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[93] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[940] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[941] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[942] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[943] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[944] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[945] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[946] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[947] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[948] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[949] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[94] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[950] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[951] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[952] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[953] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[954] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[955] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[956] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[957] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[958] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[959] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[95] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[960] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[961] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[962] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[963] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[964] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[965] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[966] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[967] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[968] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[969] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[96] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[970] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[971] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[972] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[973] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[974] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[975] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[976] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[977] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[978] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[979] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[97] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[980] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[981] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[982] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[983] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[984] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[985] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[986] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[987] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[988] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[989] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[98] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[990] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[991] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[992] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[993] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[994] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[995] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[996] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[997] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[998] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[999] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[99] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/out_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:1]\f_permutation_l_/rc ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1599:1024]\f_permutation_l_/round_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [1599:0]\f_permutation_l_/round_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \f_permutation_l_/update ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[0]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \i_reg[21]_i_reg_r_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_gate_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire i_reg_r_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire in_ready;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire is_last;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [511:0]out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1045]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1088]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1089]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1090]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1091]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1092]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1093]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1094]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1095]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1096]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1097]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1098]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1099]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1100]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1101]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1102]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1103]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1104]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1105]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1106]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1107]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1108]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1109]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1110]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1111]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1112]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1113]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1114]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1115]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1116]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1117]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1118]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1119]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1120]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1121]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1122]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1123]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1124]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1125]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1126]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1127]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1128]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1129]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1130]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1131]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1132]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1133]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1134]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1135]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1136]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1137]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1138]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1139]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1140]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1141]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1142]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1143]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1144]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1145]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1146]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1147]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1148]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1149]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1150]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1151]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1152]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1153]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1154]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1155]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1156]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1157]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1158]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1159]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1160]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1161]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1162]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1163]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1164]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1165]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1166]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1167]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1168]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1169]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1170]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1171]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1172]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1173]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1174]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1175]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1176]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1177]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1178]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1179]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1180]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1181]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1182]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1183]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1184]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1185]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1186]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1187]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1188]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1189]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1190]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1191]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1192]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1193]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1194]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1195]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1196]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1197]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1198]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1199]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1200]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1201]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1202]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1203]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1204]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1205]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1206]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1207]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1208]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1209]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1210]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1211]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1212]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1213]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1214]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1215]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1216]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1216]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1217]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1217]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1218]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1218]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1219]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1219]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1220]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1220]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1221]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1221]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1222]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1223]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1223]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1224]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1224]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1225]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1225]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1226]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1226]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1227]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1227]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1228]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1228]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1229]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1229]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1230]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1230]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1231]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1231]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1232]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1232]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1233]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1233]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1234]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1234]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1235]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1235]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1236]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1236]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1237]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1237]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1238]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1238]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1239]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1239]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1240]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1240]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1241]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1241]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1242]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1242]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1243]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1243]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1244]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1244]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1245]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1245]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1246]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1246]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1247]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1247]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1248]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1248]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1249]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1249]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1250]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1250]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1251]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1251]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1252]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1252]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1253]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1253]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1254]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1254]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1255]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1255]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1256]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1256]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1257]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1257]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1258]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1258]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1259]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1259]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1260]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1260]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1261]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1261]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1262]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1262]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1263]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1263]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1264]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1264]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1265]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1265]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1266]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1266]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1267]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1267]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1268]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1268]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1269]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1269]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1270]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1270]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1271]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1271]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1272]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1272]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1273]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1273]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1274]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1274]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1275]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1275]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1276]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1276]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1277]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1277]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1278]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1278]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1279]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1279]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1280]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1281]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1287]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[128]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1295]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[129]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[130]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1311]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[131]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[132]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[133]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1343]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1347]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[134]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[135]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[136]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[137]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[138]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[139]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1408]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1408]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1409]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1409]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[140]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1410]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1410]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1411]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1412]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1412]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1413]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1413]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1414]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1414]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1415]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1415]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1415]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1416]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1416]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1417]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1417]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1418]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1418]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1419]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1419]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[141]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1420]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1420]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1421]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1421]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1422]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1422]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1423]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1423]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1424]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1424]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1425]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1425]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1426]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1426]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1427]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1427]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1428]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1428]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1429]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1429]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[142]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1430]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1430]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1431]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1431]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1432]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1432]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1433]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1433]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1434]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1434]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1435]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1435]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1436]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1436]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1437]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1437]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1438]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1438]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1439]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1439]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[143]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1440]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1440]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1441]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1441]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1442]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1442]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1443]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1443]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1444]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1444]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1445]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1445]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1446]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1446]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1447]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1447]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1447]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1448]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1448]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1449]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1449]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[144]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1450]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1450]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1451]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1451]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1452]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1452]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1453]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1453]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1454]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1454]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1455]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1455]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1456]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1456]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1457]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1457]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1458]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1458]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1459]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1459]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[145]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1460]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1460]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1461]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1461]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1462]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1462]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1463]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1463]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1464]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1464]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1465]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1465]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1466]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1466]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1467]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1467]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1468]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1468]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1469]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1469]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[146]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1470]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1470]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1471]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1471]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1472]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1472]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1473]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1474]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1474]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1475]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1476]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1476]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1477]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1477]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1478]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1478]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1479]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[147]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1480]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1480]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1481]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1481]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1482]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1482]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1483]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1483]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1484]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1484]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1485]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1485]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1486]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1486]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1487]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1488]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1488]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1489]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1489]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[148]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1490]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1490]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1491]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1491]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1492]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1492]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1493]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1493]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1494]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1494]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1495]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1495]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1496]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1496]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1497]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1497]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1498]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1498]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1499]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1499]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[149]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1500]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1500]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1501]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1501]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1502]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1502]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1503]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1504]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1504]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1505]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1505]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1506]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1506]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1507]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1507]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1508]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1508]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1509]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1509]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[150]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1510]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1510]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1511]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1511]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1512]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1512]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1513]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1513]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1514]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1514]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1515]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1515]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1516]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1516]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1517]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1517]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1518]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1518]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1519]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1519]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[151]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1520]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1520]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1521]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1521]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1522]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1522]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1523]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1523]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1524]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1524]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1525]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1525]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1526]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1526]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1527]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1527]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1528]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1528]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1529]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1529]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[152]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1530]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1530]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1531]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1531]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1532]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1532]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1533]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1533]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1534]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1534]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1535]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1536]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1537]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1538]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1539]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[153]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1540]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1541]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1542]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1543]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1544]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1545]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1546]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1547]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1548]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1549]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[154]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1550]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1551]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1552]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1553]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1554]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1555]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1556]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1557]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1558]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1559]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[155]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1560]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1561]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1562]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1563]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1564]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1565]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1566]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1567]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1568]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1569]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[156]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1570]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1571]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1572]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1573]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1574]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1575]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1576]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1577]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1578]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1579]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[157]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1580]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1581]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1582]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1583]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1584]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1585]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1586]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1587]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1588]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1589]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[158]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1590]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1591]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1592]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1593]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1594]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1595]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1596]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1597]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1598]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[1599]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[159]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[160]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[161]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[162]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[163]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[164]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[165]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[166]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[167]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[168]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[169]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[170]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[171]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[172]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[173]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[174]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[175]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[176]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[177]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[178]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[179]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[180]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[181]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[182]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[183]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[184]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[185]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[186]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[187]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[188]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[189]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[190]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[191]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[192]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[193]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[194]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[195]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[196]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[197]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[198]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[199]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[200]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[201]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[202]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[203]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[204]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[205]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[206]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[207]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[208]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[209]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[210]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[211]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[212]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[213]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[214]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[215]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[216]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[217]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[218]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[219]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[220]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[221]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[222]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[223]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[224]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[225]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[226]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[227]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[228]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[229]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[230]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[231]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[232]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[233]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[234]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[235]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[236]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[237]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[238]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[239]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[240]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[241]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[242]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[243]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[244]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[245]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[246]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[247]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[248]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[249]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[250]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[251]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[252]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[253]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[254]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[255]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[256]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[257]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[258]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[259]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[260]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[261]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[262]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[263]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[264]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[265]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[266]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[267]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[268]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[269]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[270]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[271]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[272]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[273]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[274]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[275]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[276]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[277]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[278]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[279]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[280]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[281]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[282]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[283]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[284]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[285]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[286]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[287]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[288]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[289]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[290]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[291]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[292]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[293]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[294]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[295]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[296]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[297]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[298]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[299]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[300]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[301]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[302]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[303]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[304]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[305]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[306]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[307]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[308]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[309]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[310]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[311]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[312]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[313]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[314]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[315]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[316]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[317]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[318]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[319]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[448]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[449]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[450]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[451]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[452]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[453]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[454]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[455]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[456]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[457]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[458]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[459]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[460]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[461]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[462]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[463]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[464]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[465]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[466]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[467]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[468]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[469]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[470]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[471]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[472]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[473]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[474]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[475]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[476]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[477]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[478]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[479]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[480]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[481]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[482]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[483]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[484]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[485]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[486]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[487]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[488]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[489]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[490]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[491]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[492]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[493]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[494]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[495]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[496]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[497]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[498]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[499]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[500]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[501]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[502]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[503]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[504]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[505]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[506]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[507]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[508]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[509]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[510]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[511]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[512]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[513]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[514]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[515]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[516]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[517]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[518]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[519]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[520]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[521]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[522]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[523]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[524]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[525]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[526]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[527]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[528]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[529]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[530]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[531]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[532]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[533]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[534]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[535]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[536]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[537]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[538]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[539]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[540]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[541]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[542]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[543]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[544]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[545]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[546]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[547]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[548]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[549]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[550]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[551]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[552]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[553]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[554]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[555]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[556]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[557]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[558]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[559]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[560]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[561]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[562]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[563]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[564]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[565]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[566]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[567]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[568]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[569]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[570]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[571]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[572]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[573]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[574]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[575]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[576]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[577]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[578]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[579]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[580]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[581]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[582]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[583]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[584]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[585]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[586]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[587]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[588]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[589]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[590]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[591]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[592]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[593]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[594]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[595]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[596]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[597]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[598]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[599]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[600]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[601]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[602]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[603]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[604]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[605]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[606]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[607]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[608]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[609]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[610]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[611]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[612]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[613]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[614]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[615]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[616]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[617]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[618]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[619]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[620]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[621]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[622]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[623]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[624]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[625]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[626]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[627]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[628]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[629]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[630]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[631]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[632]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[633]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[634]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[635]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[636]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[637]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[638]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[639]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[734]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[768]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[769]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[770]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[771]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[772]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[773]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[774]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[775]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[776]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[777]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[778]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[779]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[780]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[781]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[782]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[783]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[784]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[785]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[786]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[787]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[788]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[789]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[790]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[791]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[792]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[793]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[794]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[795]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[796]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[797]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[798]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[799]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[800]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[801]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[802]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[803]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[804]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[805]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[806]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[807]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[808]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[809]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[810]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[811]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[812]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[813]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[814]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[815]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[816]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[817]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[818]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[819]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[820]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[821]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[822]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[823]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[824]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[825]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[826]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[827]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[828]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[829]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[830]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[831]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[832]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[833]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[834]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[835]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[836]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[837]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[838]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[839]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[840]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[841]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[842]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[843]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[844]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[845]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[846]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[847]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[848]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[849]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[850]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[851]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[852]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[853]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[854]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[855]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[856]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[857]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[858]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[859]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[860]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[861]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[863]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[864]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[865]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[866]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[867]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[868]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[869]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[870]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[871]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[872]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[873]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[874]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[875]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[876]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[877]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[878]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[879]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[880]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[881]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[882]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[883]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[884]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[885]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[886]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[887]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[888]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[889]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[890]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[891]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[892]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[893]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[894]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[895]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[896]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[897]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[898]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[899]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[900]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[901]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[902]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[903]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[904]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[905]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[906]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[907]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[908]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[909]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[910]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[911]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[911]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[912]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[913]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[914]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[915]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[916]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[917]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[918]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[919]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[920]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[921]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[922]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[923]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[924]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[925]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[926]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[927]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[928]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[929]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[930]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[931]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[932]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[933]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[934]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[935]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[936]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[937]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[938]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[939]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[940]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[941]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[942]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[943]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[944]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[945]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[946]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[947]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[948]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[949]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[950]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[951]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[952]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[953]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[954]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[955]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[956]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[957]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[958]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \out[959]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire out_ready;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire out_ready_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire p_0_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]p_1_out;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/done ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/i_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/out_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \padder_l_/update__1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [575:0]padder_out_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire state_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire update__0_i_1_n_0;

  assign backdoor =  update__0_i_1_n_0 ;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBA)) 
    calc_i_1
       (.I0(update__0_i_1_n_0),
        .I1(\f_permutation_l_/p_0_in ),
        .I2(\f_permutation_l_/calc ),
        .O(\f_permutation_l_/calc0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hF8)) 
    done_i_1
       (.I0(buffer_full),
        .I1(state),
        .I2(\padder_l_/done ),
        .O(done_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/calc_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/calc0 ),
        .Q(\f_permutation_l_/calc ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\i[0]_i_1__0_n_0 ),
        .Q(\f_permutation_l_/i_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[9] ),
        .Q(\f_permutation_l_/i_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[10] ),
        .Q(\f_permutation_l_/i_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[11] ),
        .Q(\f_permutation_l_/i_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[12] ),
        .Q(\f_permutation_l_/i_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[13] ),
        .Q(\f_permutation_l_/i_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[14] ),
        .Q(\f_permutation_l_/i_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[15] ),
        .Q(\f_permutation_l_/i_reg_n_0_[16] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[16] ),
        .Q(\f_permutation_l_/i_reg_n_0_[17] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[17] ),
        .Q(\f_permutation_l_/i_reg_n_0_[18] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[18] ),
        .Q(\f_permutation_l_/i_reg_n_0_[19] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_ ),
        .Q(\f_permutation_l_/i_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[19] ),
        .Q(\f_permutation_l_/i_reg_n_0_[20] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[20] ),
        .Q(\f_permutation_l_/i_reg_n_0_[21] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[21] ),
        .Q(\f_permutation_l_/p_0_in ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[1] ),
        .Q(\f_permutation_l_/i_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[2] ),
        .Q(\f_permutation_l_/i_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[3] ),
        .Q(\f_permutation_l_/i_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[4] ),
        .Q(\f_permutation_l_/i_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[5] ),
        .Q(\f_permutation_l_/i_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[6] ),
        .Q(\f_permutation_l_/i_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[7] ),
        .Q(\f_permutation_l_/i_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/i_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\f_permutation_l_/i_reg_n_0_[8] ),
        .Q(\f_permutation_l_/i_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[0] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [0]),
        .Q(\f_permutation_l_/out_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1000] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1000]),
        .Q(\f_permutation_l_/out_reg_n_0_[1000] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1001] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1001]),
        .Q(\f_permutation_l_/out_reg_n_0_[1001] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1002] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1002]),
        .Q(\f_permutation_l_/out_reg_n_0_[1002] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1003] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1003]),
        .Q(\f_permutation_l_/out_reg_n_0_[1003] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1004] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1004]),
        .Q(\f_permutation_l_/out_reg_n_0_[1004] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1005] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1005]),
        .Q(\f_permutation_l_/out_reg_n_0_[1005] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1006] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1006]),
        .Q(\f_permutation_l_/out_reg_n_0_[1006] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1007] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1007]),
        .Q(\f_permutation_l_/out_reg_n_0_[1007] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1008] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1008]),
        .Q(\f_permutation_l_/out_reg_n_0_[1008] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1009] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1009]),
        .Q(\f_permutation_l_/out_reg_n_0_[1009] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[100] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [100]),
        .Q(\f_permutation_l_/out_reg_n_0_[100] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1010] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1010]),
        .Q(\f_permutation_l_/out_reg_n_0_[1010] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1011] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1011]),
        .Q(\f_permutation_l_/out_reg_n_0_[1011] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1012] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1012]),
        .Q(\f_permutation_l_/out_reg_n_0_[1012] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1013] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1013]),
        .Q(\f_permutation_l_/out_reg_n_0_[1013] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1014] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1014]),
        .Q(\f_permutation_l_/out_reg_n_0_[1014] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1015] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1015]),
        .Q(\f_permutation_l_/out_reg_n_0_[1015] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1016] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1016]),
        .Q(\f_permutation_l_/out_reg_n_0_[1016] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1017] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1017]),
        .Q(\f_permutation_l_/out_reg_n_0_[1017] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1018] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1018]),
        .Q(\f_permutation_l_/out_reg_n_0_[1018] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1019] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1019]),
        .Q(\f_permutation_l_/out_reg_n_0_[1019] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[101] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [101]),
        .Q(\f_permutation_l_/out_reg_n_0_[101] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1020] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1020]),
        .Q(\f_permutation_l_/out_reg_n_0_[1020] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1021] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1021]),
        .Q(\f_permutation_l_/out_reg_n_0_[1021] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1022] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1022]),
        .Q(\f_permutation_l_/out_reg_n_0_[1022] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1023] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1023]),
        .Q(\f_permutation_l_/out_reg_n_0_[1023] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1024] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1024]),
        .Q(\f_permutation_l_/out_reg_n_0_[1024] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1025] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1025]),
        .Q(\f_permutation_l_/out_reg_n_0_[1025] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1026] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1026]),
        .Q(\f_permutation_l_/out_reg_n_0_[1026] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1027] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1027]),
        .Q(\f_permutation_l_/out_reg_n_0_[1027] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1028] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1028]),
        .Q(\f_permutation_l_/out_reg_n_0_[1028] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1029] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1029]),
        .Q(\f_permutation_l_/out_reg_n_0_[1029] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[102] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [102]),
        .Q(\f_permutation_l_/out_reg_n_0_[102] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1030] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1030]),
        .Q(\f_permutation_l_/out_reg_n_0_[1030] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1031] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1031]),
        .Q(\f_permutation_l_/out_reg_n_0_[1031] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1032] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1032]),
        .Q(\f_permutation_l_/out_reg_n_0_[1032] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1033] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1033]),
        .Q(\f_permutation_l_/out_reg_n_0_[1033] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1034] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1034]),
        .Q(\f_permutation_l_/out_reg_n_0_[1034] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1035] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1035]),
        .Q(\f_permutation_l_/out_reg_n_0_[1035] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1036] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1036]),
        .Q(\f_permutation_l_/out_reg_n_0_[1036] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1037] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1037]),
        .Q(\f_permutation_l_/out_reg_n_0_[1037] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1038] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1038]),
        .Q(\f_permutation_l_/out_reg_n_0_[1038] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1039] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1039]),
        .Q(\f_permutation_l_/out_reg_n_0_[1039] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[103] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [103]),
        .Q(\f_permutation_l_/out_reg_n_0_[103] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1040] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1040]),
        .Q(\f_permutation_l_/out_reg_n_0_[1040] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1041] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1041]),
        .Q(\f_permutation_l_/out_reg_n_0_[1041] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1042] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1042]),
        .Q(\f_permutation_l_/out_reg_n_0_[1042] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1043] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1043]),
        .Q(\f_permutation_l_/out_reg_n_0_[1043] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1044] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1044]),
        .Q(\f_permutation_l_/out_reg_n_0_[1044] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1045] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1045]),
        .Q(\f_permutation_l_/out_reg_n_0_[1045] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1046] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1046]),
        .Q(\f_permutation_l_/out_reg_n_0_[1046] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1047] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1047]),
        .Q(\f_permutation_l_/out_reg_n_0_[1047] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1048] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1048]),
        .Q(\f_permutation_l_/out_reg_n_0_[1048] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1049] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1049]),
        .Q(\f_permutation_l_/out_reg_n_0_[1049] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[104] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [104]),
        .Q(\f_permutation_l_/out_reg_n_0_[104] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1050] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1050]),
        .Q(\f_permutation_l_/out_reg_n_0_[1050] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1051] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1051]),
        .Q(\f_permutation_l_/out_reg_n_0_[1051] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1052] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1052]),
        .Q(\f_permutation_l_/out_reg_n_0_[1052] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1053] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1053]),
        .Q(\f_permutation_l_/out_reg_n_0_[1053] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1054] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1054]),
        .Q(\f_permutation_l_/out_reg_n_0_[1054] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1055] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1055]),
        .Q(\f_permutation_l_/out_reg_n_0_[1055] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1056] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1056]),
        .Q(\f_permutation_l_/out_reg_n_0_[1056] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1057] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1057]),
        .Q(\f_permutation_l_/out_reg_n_0_[1057] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1058] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1058]),
        .Q(\f_permutation_l_/out_reg_n_0_[1058] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1059] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1059]),
        .Q(\f_permutation_l_/out_reg_n_0_[1059] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[105] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [105]),
        .Q(\f_permutation_l_/out_reg_n_0_[105] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1060] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1060]),
        .Q(\f_permutation_l_/out_reg_n_0_[1060] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1061] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1061]),
        .Q(\f_permutation_l_/out_reg_n_0_[1061] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1062] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1062]),
        .Q(\f_permutation_l_/out_reg_n_0_[1062] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1063] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1063]),
        .Q(\f_permutation_l_/out_reg_n_0_[1063] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1064] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1064]),
        .Q(\f_permutation_l_/out_reg_n_0_[1064] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1065] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1065]),
        .Q(\f_permutation_l_/out_reg_n_0_[1065] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1066] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1066]),
        .Q(\f_permutation_l_/out_reg_n_0_[1066] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1067] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1067]),
        .Q(\f_permutation_l_/out_reg_n_0_[1067] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1068] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1068]),
        .Q(\f_permutation_l_/out_reg_n_0_[1068] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1069] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1069]),
        .Q(\f_permutation_l_/out_reg_n_0_[1069] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[106] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [106]),
        .Q(\f_permutation_l_/out_reg_n_0_[106] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1070] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1070]),
        .Q(\f_permutation_l_/out_reg_n_0_[1070] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1071] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1071]),
        .Q(\f_permutation_l_/out_reg_n_0_[1071] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1072] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1072]),
        .Q(\f_permutation_l_/out_reg_n_0_[1072] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1073] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1073]),
        .Q(\f_permutation_l_/out_reg_n_0_[1073] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1074] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1074]),
        .Q(\f_permutation_l_/out_reg_n_0_[1074] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1075] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1075]),
        .Q(\f_permutation_l_/out_reg_n_0_[1075] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1076] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1076]),
        .Q(\f_permutation_l_/out_reg_n_0_[1076] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1077] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1077]),
        .Q(\f_permutation_l_/out_reg_n_0_[1077] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1078] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1078]),
        .Q(\f_permutation_l_/out_reg_n_0_[1078] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1079] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1079]),
        .Q(\f_permutation_l_/out_reg_n_0_[1079] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[107] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [107]),
        .Q(\f_permutation_l_/out_reg_n_0_[107] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1080] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1080]),
        .Q(\f_permutation_l_/out_reg_n_0_[1080] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1081] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1081]),
        .Q(\f_permutation_l_/out_reg_n_0_[1081] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1082] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1082]),
        .Q(\f_permutation_l_/out_reg_n_0_[1082] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1083] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1083]),
        .Q(\f_permutation_l_/out_reg_n_0_[1083] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1084] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1084]),
        .Q(\f_permutation_l_/out_reg_n_0_[1084] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1085] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1085]),
        .Q(\f_permutation_l_/out_reg_n_0_[1085] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1086] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1086]),
        .Q(\f_permutation_l_/out_reg_n_0_[1086] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1087] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1087]),
        .Q(\f_permutation_l_/out_reg_n_0_[1087] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1088] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1088]),
        .Q(out[56]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1089] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1089]),
        .Q(out[57]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[108] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [108]),
        .Q(\f_permutation_l_/out_reg_n_0_[108] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1090] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1090]),
        .Q(out[58]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1091] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1091]),
        .Q(out[59]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1092] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1092]),
        .Q(out[60]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1093] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1093]),
        .Q(out[61]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1094] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1094]),
        .Q(out[62]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1095] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1095]),
        .Q(out[63]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1096] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1096]),
        .Q(out[48]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1097] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1097]),
        .Q(out[49]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1098] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1098]),
        .Q(out[50]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1099] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1099]),
        .Q(out[51]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[109] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [109]),
        .Q(\f_permutation_l_/out_reg_n_0_[109] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[10] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [10]),
        .Q(\f_permutation_l_/out_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1100] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1100]),
        .Q(out[52]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1101] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1101]),
        .Q(out[53]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1102] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1102]),
        .Q(out[54]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1103] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1103]),
        .Q(out[55]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1104] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1104]),
        .Q(out[40]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1105] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1105]),
        .Q(out[41]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1106] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1106]),
        .Q(out[42]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1107] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1107]),
        .Q(out[43]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1108] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1108]),
        .Q(out[44]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1109] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1109]),
        .Q(out[45]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[110] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [110]),
        .Q(\f_permutation_l_/out_reg_n_0_[110] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1110] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1110]),
        .Q(out[46]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1111] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1111]),
        .Q(out[47]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1112] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1112]),
        .Q(out[32]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1113] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1113]),
        .Q(out[33]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1114] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1114]),
        .Q(out[34]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1115] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1115]),
        .Q(out[35]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1116] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1116]),
        .Q(out[36]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1117] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1117]),
        .Q(out[37]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1118] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1118]),
        .Q(out[38]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1119] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1119]),
        .Q(out[39]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[111] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [111]),
        .Q(\f_permutation_l_/out_reg_n_0_[111] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1120] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1120]),
        .Q(out[24]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1121] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1121]),
        .Q(out[25]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1122] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1122]),
        .Q(out[26]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1123] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1123]),
        .Q(out[27]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1124] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1124]),
        .Q(out[28]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1125] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1125]),
        .Q(out[29]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1126] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1126]),
        .Q(out[30]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1127] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1127]),
        .Q(out[31]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1128] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1128]),
        .Q(out[16]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1129] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1129]),
        .Q(out[17]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[112] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [112]),
        .Q(\f_permutation_l_/out_reg_n_0_[112] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1130] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1130]),
        .Q(out[18]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1131] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1131]),
        .Q(out[19]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1132] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1132]),
        .Q(out[20]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1133] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1133]),
        .Q(out[21]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1134] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1134]),
        .Q(out[22]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1135] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1135]),
        .Q(out[23]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1136] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1136]),
        .Q(out[8]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1137] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1137]),
        .Q(out[9]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1138] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1138]),
        .Q(out[10]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1139] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1139]),
        .Q(out[11]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[113] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [113]),
        .Q(\f_permutation_l_/out_reg_n_0_[113] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1140] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1140]),
        .Q(out[12]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1141] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1141]),
        .Q(out[13]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1142] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1142]),
        .Q(out[14]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1143] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1143]),
        .Q(out[15]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1144] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1144]),
        .Q(out[0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1145] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1145]),
        .Q(out[1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1146] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1146]),
        .Q(out[2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1147] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1147]),
        .Q(out[3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1148] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1148]),
        .Q(out[4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1149] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1149]),
        .Q(out[5]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[114] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [114]),
        .Q(\f_permutation_l_/out_reg_n_0_[114] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1150] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1150]),
        .Q(out[6]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1151] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1151]),
        .Q(out[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1152] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1152]),
        .Q(out[120]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1153] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1153]),
        .Q(out[121]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1154] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1154]),
        .Q(out[122]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1155] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1155]),
        .Q(out[123]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1156] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1156]),
        .Q(out[124]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1157] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1157]),
        .Q(out[125]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1158] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1158]),
        .Q(out[126]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1159] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1159]),
        .Q(out[127]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[115] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [115]),
        .Q(\f_permutation_l_/out_reg_n_0_[115] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1160] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1160]),
        .Q(out[112]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1161] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1161]),
        .Q(out[113]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1162] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1162]),
        .Q(out[114]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1163] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1163]),
        .Q(out[115]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1164] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1164]),
        .Q(out[116]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1165] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1165]),
        .Q(out[117]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1166] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1166]),
        .Q(out[118]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1167] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1167]),
        .Q(out[119]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1168] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1168]),
        .Q(out[104]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1169] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1169]),
        .Q(out[105]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[116] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [116]),
        .Q(\f_permutation_l_/out_reg_n_0_[116] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1170] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1170]),
        .Q(out[106]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1171] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1171]),
        .Q(out[107]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1172] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1172]),
        .Q(out[108]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1173] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1173]),
        .Q(out[109]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1174] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1174]),
        .Q(out[110]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1175] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1175]),
        .Q(out[111]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1176] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1176]),
        .Q(out[96]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1177] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1177]),
        .Q(out[97]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1178] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1178]),
        .Q(out[98]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1179] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1179]),
        .Q(out[99]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[117] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [117]),
        .Q(\f_permutation_l_/out_reg_n_0_[117] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1180] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1180]),
        .Q(out[100]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1181] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1181]),
        .Q(out[101]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1182] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1182]),
        .Q(out[102]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1183] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1183]),
        .Q(out[103]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1184] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1184]),
        .Q(out[88]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1185] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1185]),
        .Q(out[89]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1186] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1186]),
        .Q(out[90]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1187] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1187]),
        .Q(out[91]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1188] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1188]),
        .Q(out[92]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1189] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1189]),
        .Q(out[93]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[118] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [118]),
        .Q(\f_permutation_l_/out_reg_n_0_[118] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1190] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1190]),
        .Q(out[94]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1191] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1191]),
        .Q(out[95]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1192] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1192]),
        .Q(out[80]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1193] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1193]),
        .Q(out[81]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1194] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1194]),
        .Q(out[82]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1195] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1195]),
        .Q(out[83]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1196] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1196]),
        .Q(out[84]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1197] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1197]),
        .Q(out[85]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1198] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1198]),
        .Q(out[86]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1199] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1199]),
        .Q(out[87]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[119] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [119]),
        .Q(\f_permutation_l_/out_reg_n_0_[119] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[11] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [11]),
        .Q(\f_permutation_l_/out_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1200] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1200]),
        .Q(out[72]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1201] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1201]),
        .Q(out[73]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1202] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1202]),
        .Q(out[74]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1203] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1203]),
        .Q(out[75]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1204] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1204]),
        .Q(out[76]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1205] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1205]),
        .Q(out[77]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1206] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1206]),
        .Q(out[78]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1207] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1207]),
        .Q(out[79]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1208] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1208]),
        .Q(out[64]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1209] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1209]),
        .Q(out[65]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[120] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [120]),
        .Q(\f_permutation_l_/out_reg_n_0_[120] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1210] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1210]),
        .Q(out[66]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1211] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1211]),
        .Q(out[67]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1212] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1212]),
        .Q(out[68]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1213] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1213]),
        .Q(out[69]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1214] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1214]),
        .Q(out[70]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1215] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1215]),
        .Q(out[71]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1216] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1216]),
        .Q(out[184]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1217] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1217]),
        .Q(out[185]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1218] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1218]),
        .Q(out[186]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1219] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1219]),
        .Q(out[187]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[121] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [121]),
        .Q(\f_permutation_l_/out_reg_n_0_[121] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1220] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1220]),
        .Q(out[188]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1221] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1221]),
        .Q(out[189]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1222] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1222]),
        .Q(out[190]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1223] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1223]),
        .Q(out[191]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1224] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1224]),
        .Q(out[176]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1225] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1225]),
        .Q(out[177]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1226] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1226]),
        .Q(out[178]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1227] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1227]),
        .Q(out[179]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1228] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1228]),
        .Q(out[180]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1229] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1229]),
        .Q(out[181]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[122] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [122]),
        .Q(\f_permutation_l_/out_reg_n_0_[122] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1230] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1230]),
        .Q(out[182]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1231] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1231]),
        .Q(out[183]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1232] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1232]),
        .Q(out[168]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1233] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1233]),
        .Q(out[169]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1234] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1234]),
        .Q(out[170]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1235] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1235]),
        .Q(out[171]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1236] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1236]),
        .Q(out[172]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1237] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1237]),
        .Q(out[173]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1238] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1238]),
        .Q(out[174]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1239] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1239]),
        .Q(out[175]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[123] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [123]),
        .Q(\f_permutation_l_/out_reg_n_0_[123] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1240] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1240]),
        .Q(out[160]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1241] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1241]),
        .Q(out[161]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1242] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1242]),
        .Q(out[162]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1243] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1243]),
        .Q(out[163]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1244] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1244]),
        .Q(out[164]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1245] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1245]),
        .Q(out[165]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1246] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1246]),
        .Q(out[166]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1247] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1247]),
        .Q(out[167]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1248] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1248]),
        .Q(out[152]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1249] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1249]),
        .Q(out[153]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[124] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [124]),
        .Q(\f_permutation_l_/out_reg_n_0_[124] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1250] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1250]),
        .Q(out[154]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1251] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1251]),
        .Q(out[155]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1252] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1252]),
        .Q(out[156]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1253] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1253]),
        .Q(out[157]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1254] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1254]),
        .Q(out[158]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1255] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1255]),
        .Q(out[159]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1256] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1256]),
        .Q(out[144]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1257] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1257]),
        .Q(out[145]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1258] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1258]),
        .Q(out[146]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1259] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1259]),
        .Q(out[147]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[125] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [125]),
        .Q(\f_permutation_l_/out_reg_n_0_[125] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1260] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1260]),
        .Q(out[148]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1261] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1261]),
        .Q(out[149]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1262] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1262]),
        .Q(out[150]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1263] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1263]),
        .Q(out[151]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1264] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1264]),
        .Q(out[136]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1265] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1265]),
        .Q(out[137]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1266] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1266]),
        .Q(out[138]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1267] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1267]),
        .Q(out[139]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1268] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1268]),
        .Q(out[140]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1269] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1269]),
        .Q(out[141]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[126] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [126]),
        .Q(\f_permutation_l_/out_reg_n_0_[126] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1270] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1270]),
        .Q(out[142]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1271] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1271]),
        .Q(out[143]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1272] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1272]),
        .Q(out[128]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1273] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1273]),
        .Q(out[129]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1274] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1274]),
        .Q(out[130]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1275] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1275]),
        .Q(out[131]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1276] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1276]),
        .Q(out[132]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1277] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1277]),
        .Q(out[133]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1278] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1278]),
        .Q(out[134]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1279] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1279]),
        .Q(out[135]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[127] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [127]),
        .Q(\f_permutation_l_/out_reg_n_0_[127] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1280] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1280]),
        .Q(out[248]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1281] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1281]),
        .Q(out[249]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1282] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1282]),
        .Q(out[250]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1283] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1283]),
        .Q(out[251]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1284] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1284]),
        .Q(out[252]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1285] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1285]),
        .Q(out[253]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1286] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1286]),
        .Q(out[254]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1287] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1287]),
        .Q(out[255]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1288] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1288]),
        .Q(out[240]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1289] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1289]),
        .Q(out[241]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[128] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [128]),
        .Q(\f_permutation_l_/out_reg_n_0_[128] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1290] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1290]),
        .Q(out[242]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1291] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1291]),
        .Q(out[243]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1292] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1292]),
        .Q(out[244]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1293] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1293]),
        .Q(out[245]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1294] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1294]),
        .Q(out[246]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1295] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1295]),
        .Q(out[247]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1296] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1296]),
        .Q(out[232]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1297] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1297]),
        .Q(out[233]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1298] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1298]),
        .Q(out[234]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1299] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1299]),
        .Q(out[235]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[129] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [129]),
        .Q(\f_permutation_l_/out_reg_n_0_[129] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[12] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [12]),
        .Q(\f_permutation_l_/out_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1300] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1300]),
        .Q(out[236]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1301] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1301]),
        .Q(out[237]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1302] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1302]),
        .Q(out[238]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1303] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1303]),
        .Q(out[239]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1304] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1304]),
        .Q(out[224]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1305] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1305]),
        .Q(out[225]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1306] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1306]),
        .Q(out[226]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1307] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1307]),
        .Q(out[227]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1308] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1308]),
        .Q(out[228]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1309] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1309]),
        .Q(out[229]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[130] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [130]),
        .Q(\f_permutation_l_/out_reg_n_0_[130] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1310] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1310]),
        .Q(out[230]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1311] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1311]),
        .Q(out[231]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1312] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1312]),
        .Q(out[216]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1313] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1313]),
        .Q(out[217]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1314] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1314]),
        .Q(out[218]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1315] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1315]),
        .Q(out[219]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1316] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1316]),
        .Q(out[220]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1317] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1317]),
        .Q(out[221]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1318] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1318]),
        .Q(out[222]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1319] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1319]),
        .Q(out[223]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[131] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [131]),
        .Q(\f_permutation_l_/out_reg_n_0_[131] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1320] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1320]),
        .Q(out[208]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1321] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1321]),
        .Q(out[209]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1322] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1322]),
        .Q(out[210]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1323] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1323]),
        .Q(out[211]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1324] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1324]),
        .Q(out[212]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1325] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1325]),
        .Q(out[213]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1326] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1326]),
        .Q(out[214]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1327] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1327]),
        .Q(out[215]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1328] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1328]),
        .Q(out[200]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1329] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1329]),
        .Q(out[201]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[132] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [132]),
        .Q(\f_permutation_l_/out_reg_n_0_[132] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1330] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1330]),
        .Q(out[202]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1331] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1331]),
        .Q(out[203]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1332] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1332]),
        .Q(out[204]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1333] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1333]),
        .Q(out[205]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1334] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1334]),
        .Q(out[206]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1335] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1335]),
        .Q(out[207]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1336] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1336]),
        .Q(out[192]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1337] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1337]),
        .Q(out[193]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1338] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1338]),
        .Q(out[194]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1339] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1339]),
        .Q(out[195]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[133] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [133]),
        .Q(\f_permutation_l_/out_reg_n_0_[133] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1340] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1340]),
        .Q(out[196]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1341] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1341]),
        .Q(out[197]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1342] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1342]),
        .Q(out[198]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1343] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1343]),
        .Q(out[199]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1344] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1344]),
        .Q(out[312]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1345] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1345]),
        .Q(out[313]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1346] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1346]),
        .Q(out[314]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1347] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1347]),
        .Q(out[315]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1348] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1348]),
        .Q(out[316]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1349] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1349]),
        .Q(out[317]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[134] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [134]),
        .Q(\f_permutation_l_/out_reg_n_0_[134] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1350] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1350]),
        .Q(out[318]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1351] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1351]),
        .Q(out[319]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1352] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1352]),
        .Q(out[304]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1353] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1353]),
        .Q(out[305]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1354] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1354]),
        .Q(out[306]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1355] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1355]),
        .Q(out[307]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1356] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1356]),
        .Q(out[308]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1357] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1357]),
        .Q(out[309]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1358] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1358]),
        .Q(out[310]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1359] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1359]),
        .Q(out[311]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[135] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [135]),
        .Q(\f_permutation_l_/out_reg_n_0_[135] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1360] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1360]),
        .Q(out[296]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1361] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1361]),
        .Q(out[297]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1362] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1362]),
        .Q(out[298]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1363] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1363]),
        .Q(out[299]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1364] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1364]),
        .Q(out[300]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1365] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1365]),
        .Q(out[301]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1366] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1366]),
        .Q(out[302]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1367] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1367]),
        .Q(out[303]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1368] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1368]),
        .Q(out[288]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1369] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1369]),
        .Q(out[289]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[136] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [136]),
        .Q(\f_permutation_l_/out_reg_n_0_[136] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1370] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1370]),
        .Q(out[290]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1371] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1371]),
        .Q(out[291]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1372] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1372]),
        .Q(out[292]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1373] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1373]),
        .Q(out[293]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1374] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1374]),
        .Q(out[294]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1375] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1375]),
        .Q(out[295]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1376] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1376]),
        .Q(out[280]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1377] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1377]),
        .Q(out[281]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1378] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1378]),
        .Q(out[282]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1379] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1379]),
        .Q(out[283]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[137] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [137]),
        .Q(\f_permutation_l_/out_reg_n_0_[137] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1380] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1380]),
        .Q(out[284]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1381] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1381]),
        .Q(out[285]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1382] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1382]),
        .Q(out[286]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1383] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1383]),
        .Q(out[287]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1384] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1384]),
        .Q(out[272]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1385] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1385]),
        .Q(out[273]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1386] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1386]),
        .Q(out[274]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1387] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1387]),
        .Q(out[275]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1388] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1388]),
        .Q(out[276]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1389] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1389]),
        .Q(out[277]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[138] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [138]),
        .Q(\f_permutation_l_/out_reg_n_0_[138] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1390] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1390]),
        .Q(out[278]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1391] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1391]),
        .Q(out[279]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1392] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1392]),
        .Q(out[264]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1393] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1393]),
        .Q(out[265]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1394] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1394]),
        .Q(out[266]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1395] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1395]),
        .Q(out[267]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1396] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1396]),
        .Q(out[268]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1397] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1397]),
        .Q(out[269]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1398] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1398]),
        .Q(out[270]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1399] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1399]),
        .Q(out[271]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[139] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [139]),
        .Q(\f_permutation_l_/out_reg_n_0_[139] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[13] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [13]),
        .Q(\f_permutation_l_/out_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1400] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1400]),
        .Q(out[256]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1401] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1401]),
        .Q(out[257]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1402] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1402]),
        .Q(out[258]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1403] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1403]),
        .Q(out[259]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1404] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1404]),
        .Q(out[260]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1405] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1405]),
        .Q(out[261]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1406] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1406]),
        .Q(out[262]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1407] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1407]),
        .Q(out[263]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1408] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1408]),
        .Q(out[376]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1409] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1409]),
        .Q(out[377]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[140] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [140]),
        .Q(\f_permutation_l_/out_reg_n_0_[140] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1410] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1410]),
        .Q(out[378]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1411] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1411]),
        .Q(out[379]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1412] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1412]),
        .Q(out[380]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1413] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1413]),
        .Q(out[381]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1414] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1414]),
        .Q(out[382]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1415] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1415]),
        .Q(out[383]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1416] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1416]),
        .Q(out[368]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1417] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1417]),
        .Q(out[369]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1418] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1418]),
        .Q(out[370]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1419] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1419]),
        .Q(out[371]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[141] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [141]),
        .Q(\f_permutation_l_/out_reg_n_0_[141] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1420] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1420]),
        .Q(out[372]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1421] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1421]),
        .Q(out[373]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1422] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1422]),
        .Q(out[374]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1423] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1423]),
        .Q(out[375]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1424] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1424]),
        .Q(out[360]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1425] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1425]),
        .Q(out[361]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1426] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1426]),
        .Q(out[362]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1427] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1427]),
        .Q(out[363]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1428] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1428]),
        .Q(out[364]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1429] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1429]),
        .Q(out[365]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[142] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [142]),
        .Q(\f_permutation_l_/out_reg_n_0_[142] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1430] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1430]),
        .Q(out[366]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1431] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1431]),
        .Q(out[367]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1432] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1432]),
        .Q(out[352]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1433] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1433]),
        .Q(out[353]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1434] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1434]),
        .Q(out[354]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1435] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1435]),
        .Q(out[355]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1436] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1436]),
        .Q(out[356]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1437] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1437]),
        .Q(out[357]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1438] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1438]),
        .Q(out[358]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1439] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1439]),
        .Q(out[359]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[143] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [143]),
        .Q(\f_permutation_l_/out_reg_n_0_[143] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1440] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1440]),
        .Q(out[344]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1441] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1441]),
        .Q(out[345]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1442] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1442]),
        .Q(out[346]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1443] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1443]),
        .Q(out[347]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1444] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1444]),
        .Q(out[348]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1445] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1445]),
        .Q(out[349]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1446] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1446]),
        .Q(out[350]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1447] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1447]),
        .Q(out[351]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1448] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1448]),
        .Q(out[336]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1449] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1449]),
        .Q(out[337]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[144] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [144]),
        .Q(\f_permutation_l_/out_reg_n_0_[144] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1450] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1450]),
        .Q(out[338]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1451] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1451]),
        .Q(out[339]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1452] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1452]),
        .Q(out[340]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1453] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1453]),
        .Q(out[341]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1454] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1454]),
        .Q(out[342]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1455] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1455]),
        .Q(out[343]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1456] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1456]),
        .Q(out[328]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1457] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1457]),
        .Q(out[329]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1458] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1458]),
        .Q(out[330]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1459] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1459]),
        .Q(out[331]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[145] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [145]),
        .Q(\f_permutation_l_/out_reg_n_0_[145] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1460] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1460]),
        .Q(out[332]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1461] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1461]),
        .Q(out[333]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1462] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1462]),
        .Q(out[334]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1463] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1463]),
        .Q(out[335]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1464] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1464]),
        .Q(out[320]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1465] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1465]),
        .Q(out[321]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1466] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1466]),
        .Q(out[322]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1467] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1467]),
        .Q(out[323]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1468] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1468]),
        .Q(out[324]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1469] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1469]),
        .Q(out[325]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[146] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [146]),
        .Q(\f_permutation_l_/out_reg_n_0_[146] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1470] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1470]),
        .Q(out[326]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1471] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1471]),
        .Q(out[327]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1472] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1472]),
        .Q(out[440]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1473] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1473]),
        .Q(out[441]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1474] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1474]),
        .Q(out[442]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1475] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1475]),
        .Q(out[443]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1476] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1476]),
        .Q(out[444]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1477] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1477]),
        .Q(out[445]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1478] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1478]),
        .Q(out[446]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1479] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1479]),
        .Q(out[447]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[147] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [147]),
        .Q(\f_permutation_l_/out_reg_n_0_[147] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1480] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1480]),
        .Q(out[432]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1481] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1481]),
        .Q(out[433]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1482] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1482]),
        .Q(out[434]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1483] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1483]),
        .Q(out[435]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1484] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1484]),
        .Q(out[436]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1485] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1485]),
        .Q(out[437]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1486] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1486]),
        .Q(out[438]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1487] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1487]),
        .Q(out[439]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1488] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1488]),
        .Q(out[424]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1489] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1489]),
        .Q(out[425]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[148] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [148]),
        .Q(\f_permutation_l_/out_reg_n_0_[148] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1490] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1490]),
        .Q(out[426]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1491] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1491]),
        .Q(out[427]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1492] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1492]),
        .Q(out[428]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1493] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1493]),
        .Q(out[429]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1494] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1494]),
        .Q(out[430]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1495] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1495]),
        .Q(out[431]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1496] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1496]),
        .Q(out[416]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1497] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1497]),
        .Q(out[417]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1498] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1498]),
        .Q(out[418]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1499] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1499]),
        .Q(out[419]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[149] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [149]),
        .Q(\f_permutation_l_/out_reg_n_0_[149] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[14] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [14]),
        .Q(\f_permutation_l_/out_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1500] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1500]),
        .Q(out[420]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1501] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1501]),
        .Q(out[421]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1502] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1502]),
        .Q(out[422]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1503] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1503]),
        .Q(out[423]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1504] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1504]),
        .Q(out[408]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1505] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1505]),
        .Q(out[409]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1506] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1506]),
        .Q(out[410]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1507] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1507]),
        .Q(out[411]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1508] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1508]),
        .Q(out[412]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1509] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1509]),
        .Q(out[413]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[150] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [150]),
        .Q(\f_permutation_l_/out_reg_n_0_[150] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1510] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1510]),
        .Q(out[414]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1511] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1511]),
        .Q(out[415]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1512] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1512]),
        .Q(out[400]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1513] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1513]),
        .Q(out[401]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1514] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1514]),
        .Q(out[402]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1515] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1515]),
        .Q(out[403]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1516] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1516]),
        .Q(out[404]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1517] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1517]),
        .Q(out[405]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1518] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1518]),
        .Q(out[406]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1519] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1519]),
        .Q(out[407]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[151] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [151]),
        .Q(\f_permutation_l_/out_reg_n_0_[151] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1520] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1520]),
        .Q(out[392]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1521] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1521]),
        .Q(out[393]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1522] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1522]),
        .Q(out[394]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1523] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1523]),
        .Q(out[395]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1524] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1524]),
        .Q(out[396]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1525] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1525]),
        .Q(out[397]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1526] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1526]),
        .Q(out[398]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1527] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1527]),
        .Q(out[399]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1528] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1528]),
        .Q(out[384]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1529] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1529]),
        .Q(out[385]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[152] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [152]),
        .Q(\f_permutation_l_/out_reg_n_0_[152] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1530] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1530]),
        .Q(out[386]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1531] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1531]),
        .Q(out[387]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1532] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1532]),
        .Q(out[388]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1533] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1533]),
        .Q(out[389]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1534] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1534]),
        .Q(out[390]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1535] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1535]),
        .Q(out[391]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1536] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1536]),
        .Q(out[504]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1537] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1537]),
        .Q(out[505]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1538] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1538]),
        .Q(out[506]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1539] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1539]),
        .Q(out[507]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[153] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [153]),
        .Q(\f_permutation_l_/out_reg_n_0_[153] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1540] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1540]),
        .Q(out[508]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1541] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1541]),
        .Q(out[509]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1542] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1542]),
        .Q(out[510]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1543] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1543]),
        .Q(out[511]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1544] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1544]),
        .Q(out[496]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1545] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1545]),
        .Q(out[497]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1546] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1546]),
        .Q(out[498]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1547] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1547]),
        .Q(out[499]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1548] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1548]),
        .Q(out[500]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1549] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1549]),
        .Q(out[501]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[154] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [154]),
        .Q(\f_permutation_l_/out_reg_n_0_[154] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1550] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1550]),
        .Q(out[502]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1551] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1551]),
        .Q(out[503]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1552] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1552]),
        .Q(out[488]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1553] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1553]),
        .Q(out[489]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1554] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1554]),
        .Q(out[490]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1555] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1555]),
        .Q(out[491]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1556] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1556]),
        .Q(out[492]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1557] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1557]),
        .Q(out[493]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1558] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1558]),
        .Q(out[494]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1559] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1559]),
        .Q(out[495]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[155] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [155]),
        .Q(\f_permutation_l_/out_reg_n_0_[155] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1560] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1560]),
        .Q(out[480]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1561] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1561]),
        .Q(out[481]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1562] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1562]),
        .Q(out[482]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1563] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1563]),
        .Q(out[483]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1564] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1564]),
        .Q(out[484]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1565] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1565]),
        .Q(out[485]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1566] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1566]),
        .Q(out[486]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1567] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1567]),
        .Q(out[487]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1568] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1568]),
        .Q(out[472]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1569] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1569]),
        .Q(out[473]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[156] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [156]),
        .Q(\f_permutation_l_/out_reg_n_0_[156] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1570] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1570]),
        .Q(out[474]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1571] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1571]),
        .Q(out[475]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1572] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1572]),
        .Q(out[476]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1573] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1573]),
        .Q(out[477]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1574] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1574]),
        .Q(out[478]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1575] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1575]),
        .Q(out[479]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1576] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1576]),
        .Q(out[464]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1577] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1577]),
        .Q(out[465]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1578] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1578]),
        .Q(out[466]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1579] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1579]),
        .Q(out[467]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[157] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [157]),
        .Q(\f_permutation_l_/out_reg_n_0_[157] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1580] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1580]),
        .Q(out[468]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1581] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1581]),
        .Q(out[469]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1582] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1582]),
        .Q(out[470]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1583] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1583]),
        .Q(out[471]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1584] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1584]),
        .Q(out[456]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1585] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1585]),
        .Q(out[457]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1586] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1586]),
        .Q(out[458]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1587] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1587]),
        .Q(out[459]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1588] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1588]),
        .Q(out[460]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1589] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1589]),
        .Q(out[461]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[158] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [158]),
        .Q(\f_permutation_l_/out_reg_n_0_[158] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1590] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1590]),
        .Q(out[462]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1591] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1591]),
        .Q(out[463]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1592] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1592]),
        .Q(out[448]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1593] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1593]),
        .Q(out[449]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1594] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1594]),
        .Q(out[450]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1595] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1595]),
        .Q(out[451]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1596] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1596]),
        .Q(out[452]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1597] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1597]),
        .Q(out[453]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1598] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1598]),
        .Q(out[454]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1599] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1599]),
        .Q(out[455]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[159] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [159]),
        .Q(\f_permutation_l_/out_reg_n_0_[159] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[15] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [15]),
        .Q(\f_permutation_l_/out_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[160] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [160]),
        .Q(\f_permutation_l_/out_reg_n_0_[160] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[161] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [161]),
        .Q(\f_permutation_l_/out_reg_n_0_[161] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[162] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [162]),
        .Q(\f_permutation_l_/out_reg_n_0_[162] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[163] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [163]),
        .Q(\f_permutation_l_/out_reg_n_0_[163] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[164] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [164]),
        .Q(\f_permutation_l_/out_reg_n_0_[164] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[165] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [165]),
        .Q(\f_permutation_l_/out_reg_n_0_[165] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[166] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [166]),
        .Q(\f_permutation_l_/out_reg_n_0_[166] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[167] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [167]),
        .Q(\f_permutation_l_/out_reg_n_0_[167] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[168] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [168]),
        .Q(\f_permutation_l_/out_reg_n_0_[168] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[169] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [169]),
        .Q(\f_permutation_l_/out_reg_n_0_[169] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[16] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [16]),
        .Q(\f_permutation_l_/out_reg_n_0_[16] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[170] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [170]),
        .Q(\f_permutation_l_/out_reg_n_0_[170] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[171] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [171]),
        .Q(\f_permutation_l_/out_reg_n_0_[171] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[172] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [172]),
        .Q(\f_permutation_l_/out_reg_n_0_[172] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[173] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [173]),
        .Q(\f_permutation_l_/out_reg_n_0_[173] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[174] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [174]),
        .Q(\f_permutation_l_/out_reg_n_0_[174] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[175] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [175]),
        .Q(\f_permutation_l_/out_reg_n_0_[175] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[176] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [176]),
        .Q(\f_permutation_l_/out_reg_n_0_[176] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[177] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [177]),
        .Q(\f_permutation_l_/out_reg_n_0_[177] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[178] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [178]),
        .Q(\f_permutation_l_/out_reg_n_0_[178] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[179] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [179]),
        .Q(\f_permutation_l_/out_reg_n_0_[179] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[17] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [17]),
        .Q(\f_permutation_l_/out_reg_n_0_[17] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[180] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [180]),
        .Q(\f_permutation_l_/out_reg_n_0_[180] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[181] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [181]),
        .Q(\f_permutation_l_/out_reg_n_0_[181] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[182] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [182]),
        .Q(\f_permutation_l_/out_reg_n_0_[182] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[183] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [183]),
        .Q(\f_permutation_l_/out_reg_n_0_[183] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[184] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [184]),
        .Q(\f_permutation_l_/out_reg_n_0_[184] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[185] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [185]),
        .Q(\f_permutation_l_/out_reg_n_0_[185] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[186] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [186]),
        .Q(\f_permutation_l_/out_reg_n_0_[186] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[187] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [187]),
        .Q(\f_permutation_l_/out_reg_n_0_[187] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[188] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [188]),
        .Q(\f_permutation_l_/out_reg_n_0_[188] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[189] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [189]),
        .Q(\f_permutation_l_/out_reg_n_0_[189] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[18] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [18]),
        .Q(\f_permutation_l_/out_reg_n_0_[18] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[190] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [190]),
        .Q(\f_permutation_l_/out_reg_n_0_[190] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[191] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [191]),
        .Q(\f_permutation_l_/out_reg_n_0_[191] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[192] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [192]),
        .Q(\f_permutation_l_/out_reg_n_0_[192] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[193] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [193]),
        .Q(\f_permutation_l_/out_reg_n_0_[193] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[194] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [194]),
        .Q(\f_permutation_l_/out_reg_n_0_[194] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[195] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [195]),
        .Q(\f_permutation_l_/out_reg_n_0_[195] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[196] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [196]),
        .Q(\f_permutation_l_/out_reg_n_0_[196] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[197] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [197]),
        .Q(\f_permutation_l_/out_reg_n_0_[197] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[198] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [198]),
        .Q(\f_permutation_l_/out_reg_n_0_[198] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[199] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [199]),
        .Q(\f_permutation_l_/out_reg_n_0_[199] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[19] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [19]),
        .Q(\f_permutation_l_/out_reg_n_0_[19] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[1] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [1]),
        .Q(\f_permutation_l_/out_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[200] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [200]),
        .Q(\f_permutation_l_/out_reg_n_0_[200] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[201] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [201]),
        .Q(\f_permutation_l_/out_reg_n_0_[201] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[202] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [202]),
        .Q(\f_permutation_l_/out_reg_n_0_[202] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[203] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [203]),
        .Q(\f_permutation_l_/out_reg_n_0_[203] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[204] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [204]),
        .Q(\f_permutation_l_/out_reg_n_0_[204] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[205] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [205]),
        .Q(\f_permutation_l_/out_reg_n_0_[205] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[206] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [206]),
        .Q(\f_permutation_l_/out_reg_n_0_[206] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[207] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [207]),
        .Q(\f_permutation_l_/out_reg_n_0_[207] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[208] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [208]),
        .Q(\f_permutation_l_/out_reg_n_0_[208] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[209] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [209]),
        .Q(\f_permutation_l_/out_reg_n_0_[209] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[20] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [20]),
        .Q(\f_permutation_l_/out_reg_n_0_[20] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[210] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [210]),
        .Q(\f_permutation_l_/out_reg_n_0_[210] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[211] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [211]),
        .Q(\f_permutation_l_/out_reg_n_0_[211] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[212] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [212]),
        .Q(\f_permutation_l_/out_reg_n_0_[212] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[213] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [213]),
        .Q(\f_permutation_l_/out_reg_n_0_[213] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[214] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [214]),
        .Q(\f_permutation_l_/out_reg_n_0_[214] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[215] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [215]),
        .Q(\f_permutation_l_/out_reg_n_0_[215] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[216] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [216]),
        .Q(\f_permutation_l_/out_reg_n_0_[216] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[217] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [217]),
        .Q(\f_permutation_l_/out_reg_n_0_[217] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[218] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [218]),
        .Q(\f_permutation_l_/out_reg_n_0_[218] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[219] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [219]),
        .Q(\f_permutation_l_/out_reg_n_0_[219] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[21] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [21]),
        .Q(\f_permutation_l_/out_reg_n_0_[21] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[220] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [220]),
        .Q(\f_permutation_l_/out_reg_n_0_[220] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[221] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [221]),
        .Q(\f_permutation_l_/out_reg_n_0_[221] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[222] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [222]),
        .Q(\f_permutation_l_/out_reg_n_0_[222] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[223] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [223]),
        .Q(\f_permutation_l_/out_reg_n_0_[223] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[224] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [224]),
        .Q(\f_permutation_l_/out_reg_n_0_[224] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[225] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [225]),
        .Q(\f_permutation_l_/out_reg_n_0_[225] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[226] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [226]),
        .Q(\f_permutation_l_/out_reg_n_0_[226] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[227] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [227]),
        .Q(\f_permutation_l_/out_reg_n_0_[227] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[228] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [228]),
        .Q(\f_permutation_l_/out_reg_n_0_[228] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[229] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [229]),
        .Q(\f_permutation_l_/out_reg_n_0_[229] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[22] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [22]),
        .Q(\f_permutation_l_/out_reg_n_0_[22] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[230] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [230]),
        .Q(\f_permutation_l_/out_reg_n_0_[230] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[231] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [231]),
        .Q(\f_permutation_l_/out_reg_n_0_[231] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[232] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [232]),
        .Q(\f_permutation_l_/out_reg_n_0_[232] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[233] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [233]),
        .Q(\f_permutation_l_/out_reg_n_0_[233] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[234] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [234]),
        .Q(\f_permutation_l_/out_reg_n_0_[234] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[235] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [235]),
        .Q(\f_permutation_l_/out_reg_n_0_[235] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[236] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [236]),
        .Q(\f_permutation_l_/out_reg_n_0_[236] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[237] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [237]),
        .Q(\f_permutation_l_/out_reg_n_0_[237] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[238] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [238]),
        .Q(\f_permutation_l_/out_reg_n_0_[238] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[239] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [239]),
        .Q(\f_permutation_l_/out_reg_n_0_[239] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[23] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [23]),
        .Q(\f_permutation_l_/out_reg_n_0_[23] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[240] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [240]),
        .Q(\f_permutation_l_/out_reg_n_0_[240] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[241] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [241]),
        .Q(\f_permutation_l_/out_reg_n_0_[241] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[242] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [242]),
        .Q(\f_permutation_l_/out_reg_n_0_[242] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[243] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [243]),
        .Q(\f_permutation_l_/out_reg_n_0_[243] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[244] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [244]),
        .Q(\f_permutation_l_/out_reg_n_0_[244] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[245] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [245]),
        .Q(\f_permutation_l_/out_reg_n_0_[245] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[246] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [246]),
        .Q(\f_permutation_l_/out_reg_n_0_[246] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[247] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [247]),
        .Q(\f_permutation_l_/out_reg_n_0_[247] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[248] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [248]),
        .Q(\f_permutation_l_/out_reg_n_0_[248] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[249] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [249]),
        .Q(\f_permutation_l_/out_reg_n_0_[249] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[24] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [24]),
        .Q(\f_permutation_l_/out_reg_n_0_[24] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[250] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [250]),
        .Q(\f_permutation_l_/out_reg_n_0_[250] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[251] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [251]),
        .Q(\f_permutation_l_/out_reg_n_0_[251] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[252] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [252]),
        .Q(\f_permutation_l_/out_reg_n_0_[252] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[253] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [253]),
        .Q(\f_permutation_l_/out_reg_n_0_[253] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[254] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [254]),
        .Q(\f_permutation_l_/out_reg_n_0_[254] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[255] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [255]),
        .Q(\f_permutation_l_/out_reg_n_0_[255] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[256] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [256]),
        .Q(\f_permutation_l_/out_reg_n_0_[256] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[257] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [257]),
        .Q(\f_permutation_l_/out_reg_n_0_[257] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[258] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [258]),
        .Q(\f_permutation_l_/out_reg_n_0_[258] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[259] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [259]),
        .Q(\f_permutation_l_/out_reg_n_0_[259] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[25] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [25]),
        .Q(\f_permutation_l_/out_reg_n_0_[25] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[260] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [260]),
        .Q(\f_permutation_l_/out_reg_n_0_[260] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[261] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [261]),
        .Q(\f_permutation_l_/out_reg_n_0_[261] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[262] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [262]),
        .Q(\f_permutation_l_/out_reg_n_0_[262] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[263] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [263]),
        .Q(\f_permutation_l_/out_reg_n_0_[263] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[264] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [264]),
        .Q(\f_permutation_l_/out_reg_n_0_[264] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[265] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [265]),
        .Q(\f_permutation_l_/out_reg_n_0_[265] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[266] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [266]),
        .Q(\f_permutation_l_/out_reg_n_0_[266] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[267] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [267]),
        .Q(\f_permutation_l_/out_reg_n_0_[267] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[268] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [268]),
        .Q(\f_permutation_l_/out_reg_n_0_[268] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[269] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [269]),
        .Q(\f_permutation_l_/out_reg_n_0_[269] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[26] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [26]),
        .Q(\f_permutation_l_/out_reg_n_0_[26] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[270] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [270]),
        .Q(\f_permutation_l_/out_reg_n_0_[270] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[271] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [271]),
        .Q(\f_permutation_l_/out_reg_n_0_[271] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[272] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [272]),
        .Q(\f_permutation_l_/out_reg_n_0_[272] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[273] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [273]),
        .Q(\f_permutation_l_/out_reg_n_0_[273] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[274] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [274]),
        .Q(\f_permutation_l_/out_reg_n_0_[274] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[275] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [275]),
        .Q(\f_permutation_l_/out_reg_n_0_[275] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[276] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [276]),
        .Q(\f_permutation_l_/out_reg_n_0_[276] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[277] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [277]),
        .Q(\f_permutation_l_/out_reg_n_0_[277] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[278] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [278]),
        .Q(\f_permutation_l_/out_reg_n_0_[278] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[279] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [279]),
        .Q(\f_permutation_l_/out_reg_n_0_[279] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[27] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [27]),
        .Q(\f_permutation_l_/out_reg_n_0_[27] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[280] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [280]),
        .Q(\f_permutation_l_/out_reg_n_0_[280] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[281] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [281]),
        .Q(\f_permutation_l_/out_reg_n_0_[281] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[282] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [282]),
        .Q(\f_permutation_l_/out_reg_n_0_[282] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[283] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [283]),
        .Q(\f_permutation_l_/out_reg_n_0_[283] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[284] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [284]),
        .Q(\f_permutation_l_/out_reg_n_0_[284] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[285] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [285]),
        .Q(\f_permutation_l_/out_reg_n_0_[285] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[286] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [286]),
        .Q(\f_permutation_l_/out_reg_n_0_[286] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[287] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [287]),
        .Q(\f_permutation_l_/out_reg_n_0_[287] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[288] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [288]),
        .Q(\f_permutation_l_/out_reg_n_0_[288] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[289] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [289]),
        .Q(\f_permutation_l_/out_reg_n_0_[289] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[28] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [28]),
        .Q(\f_permutation_l_/out_reg_n_0_[28] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[290] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [290]),
        .Q(\f_permutation_l_/out_reg_n_0_[290] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[291] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [291]),
        .Q(\f_permutation_l_/out_reg_n_0_[291] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[292] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [292]),
        .Q(\f_permutation_l_/out_reg_n_0_[292] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[293] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [293]),
        .Q(\f_permutation_l_/out_reg_n_0_[293] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[294] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [294]),
        .Q(\f_permutation_l_/out_reg_n_0_[294] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[295] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [295]),
        .Q(\f_permutation_l_/out_reg_n_0_[295] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[296] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [296]),
        .Q(\f_permutation_l_/out_reg_n_0_[296] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[297] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [297]),
        .Q(\f_permutation_l_/out_reg_n_0_[297] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[298] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [298]),
        .Q(\f_permutation_l_/out_reg_n_0_[298] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[299] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [299]),
        .Q(\f_permutation_l_/out_reg_n_0_[299] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[29] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [29]),
        .Q(\f_permutation_l_/out_reg_n_0_[29] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[2] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [2]),
        .Q(\f_permutation_l_/out_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[300] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [300]),
        .Q(\f_permutation_l_/out_reg_n_0_[300] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[301] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [301]),
        .Q(\f_permutation_l_/out_reg_n_0_[301] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[302] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [302]),
        .Q(\f_permutation_l_/out_reg_n_0_[302] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[303] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [303]),
        .Q(\f_permutation_l_/out_reg_n_0_[303] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[304] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [304]),
        .Q(\f_permutation_l_/out_reg_n_0_[304] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[305] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [305]),
        .Q(\f_permutation_l_/out_reg_n_0_[305] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[306] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [306]),
        .Q(\f_permutation_l_/out_reg_n_0_[306] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[307] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [307]),
        .Q(\f_permutation_l_/out_reg_n_0_[307] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[308] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [308]),
        .Q(\f_permutation_l_/out_reg_n_0_[308] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[309] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [309]),
        .Q(\f_permutation_l_/out_reg_n_0_[309] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[30] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [30]),
        .Q(\f_permutation_l_/out_reg_n_0_[30] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[310] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [310]),
        .Q(\f_permutation_l_/out_reg_n_0_[310] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[311] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [311]),
        .Q(\f_permutation_l_/out_reg_n_0_[311] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[312] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [312]),
        .Q(\f_permutation_l_/out_reg_n_0_[312] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[313] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [313]),
        .Q(\f_permutation_l_/out_reg_n_0_[313] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[314] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [314]),
        .Q(\f_permutation_l_/out_reg_n_0_[314] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[315] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [315]),
        .Q(\f_permutation_l_/out_reg_n_0_[315] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[316] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [316]),
        .Q(\f_permutation_l_/out_reg_n_0_[316] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[317] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [317]),
        .Q(\f_permutation_l_/out_reg_n_0_[317] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[318] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [318]),
        .Q(\f_permutation_l_/out_reg_n_0_[318] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[319] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [319]),
        .Q(\f_permutation_l_/out_reg_n_0_[319] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[31] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [31]),
        .Q(\f_permutation_l_/out_reg_n_0_[31] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[320] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [320]),
        .Q(\f_permutation_l_/out_reg_n_0_[320] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[321] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [321]),
        .Q(\f_permutation_l_/out_reg_n_0_[321] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[322] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [322]),
        .Q(\f_permutation_l_/out_reg_n_0_[322] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[323] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [323]),
        .Q(\f_permutation_l_/out_reg_n_0_[323] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[324] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [324]),
        .Q(\f_permutation_l_/out_reg_n_0_[324] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[325] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [325]),
        .Q(\f_permutation_l_/out_reg_n_0_[325] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[326] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [326]),
        .Q(\f_permutation_l_/out_reg_n_0_[326] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[327] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [327]),
        .Q(\f_permutation_l_/out_reg_n_0_[327] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[328] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [328]),
        .Q(\f_permutation_l_/out_reg_n_0_[328] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[329] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [329]),
        .Q(\f_permutation_l_/out_reg_n_0_[329] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[32] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [32]),
        .Q(\f_permutation_l_/out_reg_n_0_[32] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[330] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [330]),
        .Q(\f_permutation_l_/out_reg_n_0_[330] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[331] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [331]),
        .Q(\f_permutation_l_/out_reg_n_0_[331] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[332] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [332]),
        .Q(\f_permutation_l_/out_reg_n_0_[332] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[333] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [333]),
        .Q(\f_permutation_l_/out_reg_n_0_[333] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[334] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [334]),
        .Q(\f_permutation_l_/out_reg_n_0_[334] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[335] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [335]),
        .Q(\f_permutation_l_/out_reg_n_0_[335] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[336] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [336]),
        .Q(\f_permutation_l_/out_reg_n_0_[336] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[337] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [337]),
        .Q(\f_permutation_l_/out_reg_n_0_[337] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[338] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [338]),
        .Q(\f_permutation_l_/out_reg_n_0_[338] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[339] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [339]),
        .Q(\f_permutation_l_/out_reg_n_0_[339] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[33] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [33]),
        .Q(\f_permutation_l_/out_reg_n_0_[33] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[340] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [340]),
        .Q(\f_permutation_l_/out_reg_n_0_[340] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[341] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [341]),
        .Q(\f_permutation_l_/out_reg_n_0_[341] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[342] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [342]),
        .Q(\f_permutation_l_/out_reg_n_0_[342] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[343] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [343]),
        .Q(\f_permutation_l_/out_reg_n_0_[343] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[344] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [344]),
        .Q(\f_permutation_l_/out_reg_n_0_[344] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[345] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [345]),
        .Q(\f_permutation_l_/out_reg_n_0_[345] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[346] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [346]),
        .Q(\f_permutation_l_/out_reg_n_0_[346] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[347] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [347]),
        .Q(\f_permutation_l_/out_reg_n_0_[347] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[348] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [348]),
        .Q(\f_permutation_l_/out_reg_n_0_[348] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[349] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [349]),
        .Q(\f_permutation_l_/out_reg_n_0_[349] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[34] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [34]),
        .Q(\f_permutation_l_/out_reg_n_0_[34] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[350] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [350]),
        .Q(\f_permutation_l_/out_reg_n_0_[350] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[351] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [351]),
        .Q(\f_permutation_l_/out_reg_n_0_[351] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[352] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [352]),
        .Q(\f_permutation_l_/out_reg_n_0_[352] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[353] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [353]),
        .Q(\f_permutation_l_/out_reg_n_0_[353] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[354] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [354]),
        .Q(\f_permutation_l_/out_reg_n_0_[354] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[355] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [355]),
        .Q(\f_permutation_l_/out_reg_n_0_[355] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[356] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [356]),
        .Q(\f_permutation_l_/out_reg_n_0_[356] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[357] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [357]),
        .Q(\f_permutation_l_/out_reg_n_0_[357] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[358] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [358]),
        .Q(\f_permutation_l_/out_reg_n_0_[358] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[359] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [359]),
        .Q(\f_permutation_l_/out_reg_n_0_[359] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[35] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [35]),
        .Q(\f_permutation_l_/out_reg_n_0_[35] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[360] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [360]),
        .Q(\f_permutation_l_/out_reg_n_0_[360] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[361] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [361]),
        .Q(\f_permutation_l_/out_reg_n_0_[361] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[362] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [362]),
        .Q(\f_permutation_l_/out_reg_n_0_[362] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[363] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [363]),
        .Q(\f_permutation_l_/out_reg_n_0_[363] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[364] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [364]),
        .Q(\f_permutation_l_/out_reg_n_0_[364] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[365] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [365]),
        .Q(\f_permutation_l_/out_reg_n_0_[365] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[366] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [366]),
        .Q(\f_permutation_l_/out_reg_n_0_[366] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[367] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [367]),
        .Q(\f_permutation_l_/out_reg_n_0_[367] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[368] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [368]),
        .Q(\f_permutation_l_/out_reg_n_0_[368] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[369] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [369]),
        .Q(\f_permutation_l_/out_reg_n_0_[369] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[36] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [36]),
        .Q(\f_permutation_l_/out_reg_n_0_[36] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[370] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [370]),
        .Q(\f_permutation_l_/out_reg_n_0_[370] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[371] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [371]),
        .Q(\f_permutation_l_/out_reg_n_0_[371] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[372] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [372]),
        .Q(\f_permutation_l_/out_reg_n_0_[372] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[373] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [373]),
        .Q(\f_permutation_l_/out_reg_n_0_[373] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[374] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [374]),
        .Q(\f_permutation_l_/out_reg_n_0_[374] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[375] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [375]),
        .Q(\f_permutation_l_/out_reg_n_0_[375] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[376] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [376]),
        .Q(\f_permutation_l_/out_reg_n_0_[376] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[377] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [377]),
        .Q(\f_permutation_l_/out_reg_n_0_[377] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[378] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [378]),
        .Q(\f_permutation_l_/out_reg_n_0_[378] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[379] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [379]),
        .Q(\f_permutation_l_/out_reg_n_0_[379] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[37] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [37]),
        .Q(\f_permutation_l_/out_reg_n_0_[37] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[380] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [380]),
        .Q(\f_permutation_l_/out_reg_n_0_[380] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[381] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [381]),
        .Q(\f_permutation_l_/out_reg_n_0_[381] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[382] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [382]),
        .Q(\f_permutation_l_/out_reg_n_0_[382] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[383] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [383]),
        .Q(\f_permutation_l_/out_reg_n_0_[383] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[384] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [384]),
        .Q(\f_permutation_l_/out_reg_n_0_[384] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[385] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [385]),
        .Q(\f_permutation_l_/out_reg_n_0_[385] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[386] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [386]),
        .Q(\f_permutation_l_/out_reg_n_0_[386] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[387] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [387]),
        .Q(\f_permutation_l_/out_reg_n_0_[387] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[388] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [388]),
        .Q(\f_permutation_l_/out_reg_n_0_[388] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[389] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [389]),
        .Q(\f_permutation_l_/out_reg_n_0_[389] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[38] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [38]),
        .Q(\f_permutation_l_/out_reg_n_0_[38] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[390] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [390]),
        .Q(\f_permutation_l_/out_reg_n_0_[390] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[391] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [391]),
        .Q(\f_permutation_l_/out_reg_n_0_[391] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[392] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [392]),
        .Q(\f_permutation_l_/out_reg_n_0_[392] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[393] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [393]),
        .Q(\f_permutation_l_/out_reg_n_0_[393] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[394] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [394]),
        .Q(\f_permutation_l_/out_reg_n_0_[394] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[395] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [395]),
        .Q(\f_permutation_l_/out_reg_n_0_[395] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[396] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [396]),
        .Q(\f_permutation_l_/out_reg_n_0_[396] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[397] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [397]),
        .Q(\f_permutation_l_/out_reg_n_0_[397] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[398] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [398]),
        .Q(\f_permutation_l_/out_reg_n_0_[398] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[399] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [399]),
        .Q(\f_permutation_l_/out_reg_n_0_[399] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[39] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [39]),
        .Q(\f_permutation_l_/out_reg_n_0_[39] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[3] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [3]),
        .Q(\f_permutation_l_/out_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[400] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [400]),
        .Q(\f_permutation_l_/out_reg_n_0_[400] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[401] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [401]),
        .Q(\f_permutation_l_/out_reg_n_0_[401] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[402] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [402]),
        .Q(\f_permutation_l_/out_reg_n_0_[402] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[403] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [403]),
        .Q(\f_permutation_l_/out_reg_n_0_[403] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[404] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [404]),
        .Q(\f_permutation_l_/out_reg_n_0_[404] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[405] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [405]),
        .Q(\f_permutation_l_/out_reg_n_0_[405] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[406] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [406]),
        .Q(\f_permutation_l_/out_reg_n_0_[406] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[407] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [407]),
        .Q(\f_permutation_l_/out_reg_n_0_[407] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[408] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [408]),
        .Q(\f_permutation_l_/out_reg_n_0_[408] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[409] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [409]),
        .Q(\f_permutation_l_/out_reg_n_0_[409] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[40] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [40]),
        .Q(\f_permutation_l_/out_reg_n_0_[40] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[410] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [410]),
        .Q(\f_permutation_l_/out_reg_n_0_[410] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[411] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [411]),
        .Q(\f_permutation_l_/out_reg_n_0_[411] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[412] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [412]),
        .Q(\f_permutation_l_/out_reg_n_0_[412] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[413] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [413]),
        .Q(\f_permutation_l_/out_reg_n_0_[413] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[414] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [414]),
        .Q(\f_permutation_l_/out_reg_n_0_[414] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[415] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [415]),
        .Q(\f_permutation_l_/out_reg_n_0_[415] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[416] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [416]),
        .Q(\f_permutation_l_/out_reg_n_0_[416] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[417] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [417]),
        .Q(\f_permutation_l_/out_reg_n_0_[417] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[418] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [418]),
        .Q(\f_permutation_l_/out_reg_n_0_[418] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[419] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [419]),
        .Q(\f_permutation_l_/out_reg_n_0_[419] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[41] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [41]),
        .Q(\f_permutation_l_/out_reg_n_0_[41] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[420] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [420]),
        .Q(\f_permutation_l_/out_reg_n_0_[420] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[421] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [421]),
        .Q(\f_permutation_l_/out_reg_n_0_[421] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[422] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [422]),
        .Q(\f_permutation_l_/out_reg_n_0_[422] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[423] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [423]),
        .Q(\f_permutation_l_/out_reg_n_0_[423] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[424] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [424]),
        .Q(\f_permutation_l_/out_reg_n_0_[424] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[425] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [425]),
        .Q(\f_permutation_l_/out_reg_n_0_[425] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[426] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [426]),
        .Q(\f_permutation_l_/out_reg_n_0_[426] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[427] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [427]),
        .Q(\f_permutation_l_/out_reg_n_0_[427] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[428] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [428]),
        .Q(\f_permutation_l_/out_reg_n_0_[428] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[429] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [429]),
        .Q(\f_permutation_l_/out_reg_n_0_[429] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[42] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [42]),
        .Q(\f_permutation_l_/out_reg_n_0_[42] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[430] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [430]),
        .Q(\f_permutation_l_/out_reg_n_0_[430] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[431] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [431]),
        .Q(\f_permutation_l_/out_reg_n_0_[431] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[432] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [432]),
        .Q(\f_permutation_l_/out_reg_n_0_[432] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[433] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [433]),
        .Q(\f_permutation_l_/out_reg_n_0_[433] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[434] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [434]),
        .Q(\f_permutation_l_/out_reg_n_0_[434] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[435] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [435]),
        .Q(\f_permutation_l_/out_reg_n_0_[435] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[436] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [436]),
        .Q(\f_permutation_l_/out_reg_n_0_[436] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[437] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [437]),
        .Q(\f_permutation_l_/out_reg_n_0_[437] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[438] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [438]),
        .Q(\f_permutation_l_/out_reg_n_0_[438] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[439] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [439]),
        .Q(\f_permutation_l_/out_reg_n_0_[439] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[43] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [43]),
        .Q(\f_permutation_l_/out_reg_n_0_[43] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[440] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [440]),
        .Q(\f_permutation_l_/out_reg_n_0_[440] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[441] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [441]),
        .Q(\f_permutation_l_/out_reg_n_0_[441] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[442] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [442]),
        .Q(\f_permutation_l_/out_reg_n_0_[442] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[443] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [443]),
        .Q(\f_permutation_l_/out_reg_n_0_[443] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[444] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [444]),
        .Q(\f_permutation_l_/out_reg_n_0_[444] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[445] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [445]),
        .Q(\f_permutation_l_/out_reg_n_0_[445] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[446] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [446]),
        .Q(\f_permutation_l_/out_reg_n_0_[446] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[447] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [447]),
        .Q(\f_permutation_l_/out_reg_n_0_[447] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[448] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [448]),
        .Q(\f_permutation_l_/out_reg_n_0_[448] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[449] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [449]),
        .Q(\f_permutation_l_/out_reg_n_0_[449] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[44] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [44]),
        .Q(\f_permutation_l_/out_reg_n_0_[44] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[450] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [450]),
        .Q(\f_permutation_l_/out_reg_n_0_[450] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[451] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [451]),
        .Q(\f_permutation_l_/out_reg_n_0_[451] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[452] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [452]),
        .Q(\f_permutation_l_/out_reg_n_0_[452] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[453] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [453]),
        .Q(\f_permutation_l_/out_reg_n_0_[453] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[454] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [454]),
        .Q(\f_permutation_l_/out_reg_n_0_[454] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[455] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [455]),
        .Q(\f_permutation_l_/out_reg_n_0_[455] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[456] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [456]),
        .Q(\f_permutation_l_/out_reg_n_0_[456] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[457] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [457]),
        .Q(\f_permutation_l_/out_reg_n_0_[457] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[458] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [458]),
        .Q(\f_permutation_l_/out_reg_n_0_[458] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[459] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [459]),
        .Q(\f_permutation_l_/out_reg_n_0_[459] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[45] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [45]),
        .Q(\f_permutation_l_/out_reg_n_0_[45] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[460] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [460]),
        .Q(\f_permutation_l_/out_reg_n_0_[460] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[461] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [461]),
        .Q(\f_permutation_l_/out_reg_n_0_[461] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[462] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [462]),
        .Q(\f_permutation_l_/out_reg_n_0_[462] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[463] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [463]),
        .Q(\f_permutation_l_/out_reg_n_0_[463] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[464] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [464]),
        .Q(\f_permutation_l_/out_reg_n_0_[464] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[465] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [465]),
        .Q(\f_permutation_l_/out_reg_n_0_[465] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[466] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [466]),
        .Q(\f_permutation_l_/out_reg_n_0_[466] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[467] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [467]),
        .Q(\f_permutation_l_/out_reg_n_0_[467] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[468] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [468]),
        .Q(\f_permutation_l_/out_reg_n_0_[468] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[469] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [469]),
        .Q(\f_permutation_l_/out_reg_n_0_[469] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[46] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [46]),
        .Q(\f_permutation_l_/out_reg_n_0_[46] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[470] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [470]),
        .Q(\f_permutation_l_/out_reg_n_0_[470] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[471] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [471]),
        .Q(\f_permutation_l_/out_reg_n_0_[471] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[472] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [472]),
        .Q(\f_permutation_l_/out_reg_n_0_[472] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[473] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [473]),
        .Q(\f_permutation_l_/out_reg_n_0_[473] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[474] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [474]),
        .Q(\f_permutation_l_/out_reg_n_0_[474] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[475] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [475]),
        .Q(\f_permutation_l_/out_reg_n_0_[475] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[476] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [476]),
        .Q(\f_permutation_l_/out_reg_n_0_[476] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[477] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [477]),
        .Q(\f_permutation_l_/out_reg_n_0_[477] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[478] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [478]),
        .Q(\f_permutation_l_/out_reg_n_0_[478] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[479] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [479]),
        .Q(\f_permutation_l_/out_reg_n_0_[479] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[47] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [47]),
        .Q(\f_permutation_l_/out_reg_n_0_[47] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[480] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [480]),
        .Q(\f_permutation_l_/out_reg_n_0_[480] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[481] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [481]),
        .Q(\f_permutation_l_/out_reg_n_0_[481] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[482] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [482]),
        .Q(\f_permutation_l_/out_reg_n_0_[482] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[483] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [483]),
        .Q(\f_permutation_l_/out_reg_n_0_[483] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[484] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [484]),
        .Q(\f_permutation_l_/out_reg_n_0_[484] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[485] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [485]),
        .Q(\f_permutation_l_/out_reg_n_0_[485] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[486] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [486]),
        .Q(\f_permutation_l_/out_reg_n_0_[486] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[487] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [487]),
        .Q(\f_permutation_l_/out_reg_n_0_[487] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[488] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [488]),
        .Q(\f_permutation_l_/out_reg_n_0_[488] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[489] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [489]),
        .Q(\f_permutation_l_/out_reg_n_0_[489] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[48] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [48]),
        .Q(\f_permutation_l_/out_reg_n_0_[48] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[490] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [490]),
        .Q(\f_permutation_l_/out_reg_n_0_[490] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[491] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [491]),
        .Q(\f_permutation_l_/out_reg_n_0_[491] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[492] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [492]),
        .Q(\f_permutation_l_/out_reg_n_0_[492] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[493] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [493]),
        .Q(\f_permutation_l_/out_reg_n_0_[493] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[494] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [494]),
        .Q(\f_permutation_l_/out_reg_n_0_[494] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[495] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [495]),
        .Q(\f_permutation_l_/out_reg_n_0_[495] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[496] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [496]),
        .Q(\f_permutation_l_/out_reg_n_0_[496] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[497] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [497]),
        .Q(\f_permutation_l_/out_reg_n_0_[497] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[498] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [498]),
        .Q(\f_permutation_l_/out_reg_n_0_[498] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[499] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [499]),
        .Q(\f_permutation_l_/out_reg_n_0_[499] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[49] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [49]),
        .Q(\f_permutation_l_/out_reg_n_0_[49] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[4] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [4]),
        .Q(\f_permutation_l_/out_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[500] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [500]),
        .Q(\f_permutation_l_/out_reg_n_0_[500] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[501] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [501]),
        .Q(\f_permutation_l_/out_reg_n_0_[501] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[502] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [502]),
        .Q(\f_permutation_l_/out_reg_n_0_[502] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[503] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [503]),
        .Q(\f_permutation_l_/out_reg_n_0_[503] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[504] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [504]),
        .Q(\f_permutation_l_/out_reg_n_0_[504] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[505] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [505]),
        .Q(\f_permutation_l_/out_reg_n_0_[505] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[506] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [506]),
        .Q(\f_permutation_l_/out_reg_n_0_[506] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[507] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [507]),
        .Q(\f_permutation_l_/out_reg_n_0_[507] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[508] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [508]),
        .Q(\f_permutation_l_/out_reg_n_0_[508] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[509] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [509]),
        .Q(\f_permutation_l_/out_reg_n_0_[509] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[50] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [50]),
        .Q(\f_permutation_l_/out_reg_n_0_[50] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[510] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [510]),
        .Q(\f_permutation_l_/out_reg_n_0_[510] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[511] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [511]),
        .Q(\f_permutation_l_/out_reg_n_0_[511] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[512] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [512]),
        .Q(\f_permutation_l_/out_reg_n_0_[512] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[513] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [513]),
        .Q(\f_permutation_l_/out_reg_n_0_[513] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[514] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [514]),
        .Q(\f_permutation_l_/out_reg_n_0_[514] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[515] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [515]),
        .Q(\f_permutation_l_/out_reg_n_0_[515] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[516] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [516]),
        .Q(\f_permutation_l_/out_reg_n_0_[516] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[517] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [517]),
        .Q(\f_permutation_l_/out_reg_n_0_[517] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[518] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [518]),
        .Q(\f_permutation_l_/out_reg_n_0_[518] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[519] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [519]),
        .Q(\f_permutation_l_/out_reg_n_0_[519] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[51] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [51]),
        .Q(\f_permutation_l_/out_reg_n_0_[51] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[520] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [520]),
        .Q(\f_permutation_l_/out_reg_n_0_[520] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[521] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [521]),
        .Q(\f_permutation_l_/out_reg_n_0_[521] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[522] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [522]),
        .Q(\f_permutation_l_/out_reg_n_0_[522] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[523] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [523]),
        .Q(\f_permutation_l_/out_reg_n_0_[523] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[524] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [524]),
        .Q(\f_permutation_l_/out_reg_n_0_[524] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[525] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [525]),
        .Q(\f_permutation_l_/out_reg_n_0_[525] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[526] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [526]),
        .Q(\f_permutation_l_/out_reg_n_0_[526] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[527] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [527]),
        .Q(\f_permutation_l_/out_reg_n_0_[527] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[528] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [528]),
        .Q(\f_permutation_l_/out_reg_n_0_[528] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[529] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [529]),
        .Q(\f_permutation_l_/out_reg_n_0_[529] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[52] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [52]),
        .Q(\f_permutation_l_/out_reg_n_0_[52] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[530] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [530]),
        .Q(\f_permutation_l_/out_reg_n_0_[530] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[531] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [531]),
        .Q(\f_permutation_l_/out_reg_n_0_[531] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[532] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [532]),
        .Q(\f_permutation_l_/out_reg_n_0_[532] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[533] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [533]),
        .Q(\f_permutation_l_/out_reg_n_0_[533] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[534] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [534]),
        .Q(\f_permutation_l_/out_reg_n_0_[534] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[535] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [535]),
        .Q(\f_permutation_l_/out_reg_n_0_[535] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[536] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [536]),
        .Q(\f_permutation_l_/out_reg_n_0_[536] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[537] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [537]),
        .Q(\f_permutation_l_/out_reg_n_0_[537] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[538] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [538]),
        .Q(\f_permutation_l_/out_reg_n_0_[538] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[539] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [539]),
        .Q(\f_permutation_l_/out_reg_n_0_[539] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[53] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [53]),
        .Q(\f_permutation_l_/out_reg_n_0_[53] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[540] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [540]),
        .Q(\f_permutation_l_/out_reg_n_0_[540] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[541] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [541]),
        .Q(\f_permutation_l_/out_reg_n_0_[541] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[542] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [542]),
        .Q(\f_permutation_l_/out_reg_n_0_[542] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[543] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [543]),
        .Q(\f_permutation_l_/out_reg_n_0_[543] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[544] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [544]),
        .Q(\f_permutation_l_/out_reg_n_0_[544] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[545] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [545]),
        .Q(\f_permutation_l_/out_reg_n_0_[545] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[546] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [546]),
        .Q(\f_permutation_l_/out_reg_n_0_[546] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[547] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [547]),
        .Q(\f_permutation_l_/out_reg_n_0_[547] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[548] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [548]),
        .Q(\f_permutation_l_/out_reg_n_0_[548] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[549] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [549]),
        .Q(\f_permutation_l_/out_reg_n_0_[549] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[54] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [54]),
        .Q(\f_permutation_l_/out_reg_n_0_[54] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[550] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [550]),
        .Q(\f_permutation_l_/out_reg_n_0_[550] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[551] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [551]),
        .Q(\f_permutation_l_/out_reg_n_0_[551] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[552] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [552]),
        .Q(\f_permutation_l_/out_reg_n_0_[552] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[553] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [553]),
        .Q(\f_permutation_l_/out_reg_n_0_[553] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[554] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [554]),
        .Q(\f_permutation_l_/out_reg_n_0_[554] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[555] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [555]),
        .Q(\f_permutation_l_/out_reg_n_0_[555] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[556] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [556]),
        .Q(\f_permutation_l_/out_reg_n_0_[556] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[557] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [557]),
        .Q(\f_permutation_l_/out_reg_n_0_[557] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[558] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [558]),
        .Q(\f_permutation_l_/out_reg_n_0_[558] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[559] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [559]),
        .Q(\f_permutation_l_/out_reg_n_0_[559] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[55] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [55]),
        .Q(\f_permutation_l_/out_reg_n_0_[55] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[560] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [560]),
        .Q(\f_permutation_l_/out_reg_n_0_[560] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[561] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [561]),
        .Q(\f_permutation_l_/out_reg_n_0_[561] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[562] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [562]),
        .Q(\f_permutation_l_/out_reg_n_0_[562] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[563] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [563]),
        .Q(\f_permutation_l_/out_reg_n_0_[563] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[564] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [564]),
        .Q(\f_permutation_l_/out_reg_n_0_[564] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[565] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [565]),
        .Q(\f_permutation_l_/out_reg_n_0_[565] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[566] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [566]),
        .Q(\f_permutation_l_/out_reg_n_0_[566] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[567] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [567]),
        .Q(\f_permutation_l_/out_reg_n_0_[567] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[568] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [568]),
        .Q(\f_permutation_l_/out_reg_n_0_[568] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[569] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [569]),
        .Q(\f_permutation_l_/out_reg_n_0_[569] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[56] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [56]),
        .Q(\f_permutation_l_/out_reg_n_0_[56] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[570] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [570]),
        .Q(\f_permutation_l_/out_reg_n_0_[570] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[571] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [571]),
        .Q(\f_permutation_l_/out_reg_n_0_[571] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[572] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [572]),
        .Q(\f_permutation_l_/out_reg_n_0_[572] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[573] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [573]),
        .Q(\f_permutation_l_/out_reg_n_0_[573] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[574] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [574]),
        .Q(\f_permutation_l_/out_reg_n_0_[574] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[575] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [575]),
        .Q(\f_permutation_l_/out_reg_n_0_[575] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[576] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [576]),
        .Q(\f_permutation_l_/out_reg_n_0_[576] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[577] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [577]),
        .Q(\f_permutation_l_/out_reg_n_0_[577] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[578] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [578]),
        .Q(\f_permutation_l_/out_reg_n_0_[578] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[579] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [579]),
        .Q(\f_permutation_l_/out_reg_n_0_[579] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[57] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [57]),
        .Q(\f_permutation_l_/out_reg_n_0_[57] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[580] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [580]),
        .Q(\f_permutation_l_/out_reg_n_0_[580] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[581] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [581]),
        .Q(\f_permutation_l_/out_reg_n_0_[581] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[582] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [582]),
        .Q(\f_permutation_l_/out_reg_n_0_[582] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[583] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [583]),
        .Q(\f_permutation_l_/out_reg_n_0_[583] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[584] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [584]),
        .Q(\f_permutation_l_/out_reg_n_0_[584] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[585] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [585]),
        .Q(\f_permutation_l_/out_reg_n_0_[585] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[586] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [586]),
        .Q(\f_permutation_l_/out_reg_n_0_[586] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[587] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [587]),
        .Q(\f_permutation_l_/out_reg_n_0_[587] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[588] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [588]),
        .Q(\f_permutation_l_/out_reg_n_0_[588] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[589] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [589]),
        .Q(\f_permutation_l_/out_reg_n_0_[589] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[58] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [58]),
        .Q(\f_permutation_l_/out_reg_n_0_[58] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[590] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [590]),
        .Q(\f_permutation_l_/out_reg_n_0_[590] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[591] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [591]),
        .Q(\f_permutation_l_/out_reg_n_0_[591] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[592] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [592]),
        .Q(\f_permutation_l_/out_reg_n_0_[592] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[593] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [593]),
        .Q(\f_permutation_l_/out_reg_n_0_[593] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[594] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [594]),
        .Q(\f_permutation_l_/out_reg_n_0_[594] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[595] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [595]),
        .Q(\f_permutation_l_/out_reg_n_0_[595] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[596] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [596]),
        .Q(\f_permutation_l_/out_reg_n_0_[596] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[597] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [597]),
        .Q(\f_permutation_l_/out_reg_n_0_[597] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[598] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [598]),
        .Q(\f_permutation_l_/out_reg_n_0_[598] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[599] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [599]),
        .Q(\f_permutation_l_/out_reg_n_0_[599] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[59] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [59]),
        .Q(\f_permutation_l_/out_reg_n_0_[59] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[5] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [5]),
        .Q(\f_permutation_l_/out_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[600] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [600]),
        .Q(\f_permutation_l_/out_reg_n_0_[600] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[601] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [601]),
        .Q(\f_permutation_l_/out_reg_n_0_[601] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[602] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [602]),
        .Q(\f_permutation_l_/out_reg_n_0_[602] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[603] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [603]),
        .Q(\f_permutation_l_/out_reg_n_0_[603] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[604] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [604]),
        .Q(\f_permutation_l_/out_reg_n_0_[604] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[605] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [605]),
        .Q(\f_permutation_l_/out_reg_n_0_[605] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[606] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [606]),
        .Q(\f_permutation_l_/out_reg_n_0_[606] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[607] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [607]),
        .Q(\f_permutation_l_/out_reg_n_0_[607] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[608] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [608]),
        .Q(\f_permutation_l_/out_reg_n_0_[608] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[609] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [609]),
        .Q(\f_permutation_l_/out_reg_n_0_[609] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[60] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [60]),
        .Q(\f_permutation_l_/out_reg_n_0_[60] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[610] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [610]),
        .Q(\f_permutation_l_/out_reg_n_0_[610] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[611] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [611]),
        .Q(\f_permutation_l_/out_reg_n_0_[611] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[612] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [612]),
        .Q(\f_permutation_l_/out_reg_n_0_[612] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[613] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [613]),
        .Q(\f_permutation_l_/out_reg_n_0_[613] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[614] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [614]),
        .Q(\f_permutation_l_/out_reg_n_0_[614] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[615] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [615]),
        .Q(\f_permutation_l_/out_reg_n_0_[615] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[616] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [616]),
        .Q(\f_permutation_l_/out_reg_n_0_[616] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[617] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [617]),
        .Q(\f_permutation_l_/out_reg_n_0_[617] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[618] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [618]),
        .Q(\f_permutation_l_/out_reg_n_0_[618] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[619] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [619]),
        .Q(\f_permutation_l_/out_reg_n_0_[619] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[61] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [61]),
        .Q(\f_permutation_l_/out_reg_n_0_[61] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[620] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [620]),
        .Q(\f_permutation_l_/out_reg_n_0_[620] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[621] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [621]),
        .Q(\f_permutation_l_/out_reg_n_0_[621] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[622] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [622]),
        .Q(\f_permutation_l_/out_reg_n_0_[622] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[623] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [623]),
        .Q(\f_permutation_l_/out_reg_n_0_[623] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[624] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [624]),
        .Q(\f_permutation_l_/out_reg_n_0_[624] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[625] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [625]),
        .Q(\f_permutation_l_/out_reg_n_0_[625] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[626] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [626]),
        .Q(\f_permutation_l_/out_reg_n_0_[626] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[627] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [627]),
        .Q(\f_permutation_l_/out_reg_n_0_[627] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[628] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [628]),
        .Q(\f_permutation_l_/out_reg_n_0_[628] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[629] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [629]),
        .Q(\f_permutation_l_/out_reg_n_0_[629] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[62] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [62]),
        .Q(\f_permutation_l_/out_reg_n_0_[62] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[630] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [630]),
        .Q(\f_permutation_l_/out_reg_n_0_[630] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[631] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [631]),
        .Q(\f_permutation_l_/out_reg_n_0_[631] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[632] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [632]),
        .Q(\f_permutation_l_/out_reg_n_0_[632] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[633] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [633]),
        .Q(\f_permutation_l_/out_reg_n_0_[633] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[634] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [634]),
        .Q(\f_permutation_l_/out_reg_n_0_[634] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[635] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [635]),
        .Q(\f_permutation_l_/out_reg_n_0_[635] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[636] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [636]),
        .Q(\f_permutation_l_/out_reg_n_0_[636] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[637] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [637]),
        .Q(\f_permutation_l_/out_reg_n_0_[637] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[638] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [638]),
        .Q(\f_permutation_l_/out_reg_n_0_[638] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[639] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [639]),
        .Q(\f_permutation_l_/out_reg_n_0_[639] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[63] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [63]),
        .Q(\f_permutation_l_/out_reg_n_0_[63] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[640] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [640]),
        .Q(\f_permutation_l_/out_reg_n_0_[640] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[641] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [641]),
        .Q(\f_permutation_l_/out_reg_n_0_[641] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[642] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [642]),
        .Q(\f_permutation_l_/out_reg_n_0_[642] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[643] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [643]),
        .Q(\f_permutation_l_/out_reg_n_0_[643] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[644] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [644]),
        .Q(\f_permutation_l_/out_reg_n_0_[644] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[645] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [645]),
        .Q(\f_permutation_l_/out_reg_n_0_[645] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[646] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [646]),
        .Q(\f_permutation_l_/out_reg_n_0_[646] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[647] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [647]),
        .Q(\f_permutation_l_/out_reg_n_0_[647] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[648] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [648]),
        .Q(\f_permutation_l_/out_reg_n_0_[648] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[649] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [649]),
        .Q(\f_permutation_l_/out_reg_n_0_[649] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[64] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [64]),
        .Q(\f_permutation_l_/out_reg_n_0_[64] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[650] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [650]),
        .Q(\f_permutation_l_/out_reg_n_0_[650] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[651] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [651]),
        .Q(\f_permutation_l_/out_reg_n_0_[651] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[652] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [652]),
        .Q(\f_permutation_l_/out_reg_n_0_[652] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[653] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [653]),
        .Q(\f_permutation_l_/out_reg_n_0_[653] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[654] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [654]),
        .Q(\f_permutation_l_/out_reg_n_0_[654] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[655] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [655]),
        .Q(\f_permutation_l_/out_reg_n_0_[655] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[656] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [656]),
        .Q(\f_permutation_l_/out_reg_n_0_[656] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[657] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [657]),
        .Q(\f_permutation_l_/out_reg_n_0_[657] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[658] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [658]),
        .Q(\f_permutation_l_/out_reg_n_0_[658] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[659] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [659]),
        .Q(\f_permutation_l_/out_reg_n_0_[659] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[65] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [65]),
        .Q(\f_permutation_l_/out_reg_n_0_[65] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[660] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [660]),
        .Q(\f_permutation_l_/out_reg_n_0_[660] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[661] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [661]),
        .Q(\f_permutation_l_/out_reg_n_0_[661] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[662] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [662]),
        .Q(\f_permutation_l_/out_reg_n_0_[662] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[663] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [663]),
        .Q(\f_permutation_l_/out_reg_n_0_[663] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[664] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [664]),
        .Q(\f_permutation_l_/out_reg_n_0_[664] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[665] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [665]),
        .Q(\f_permutation_l_/out_reg_n_0_[665] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[666] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [666]),
        .Q(\f_permutation_l_/out_reg_n_0_[666] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[667] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [667]),
        .Q(\f_permutation_l_/out_reg_n_0_[667] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[668] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [668]),
        .Q(\f_permutation_l_/out_reg_n_0_[668] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[669] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [669]),
        .Q(\f_permutation_l_/out_reg_n_0_[669] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[66] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [66]),
        .Q(\f_permutation_l_/out_reg_n_0_[66] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[670] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [670]),
        .Q(\f_permutation_l_/out_reg_n_0_[670] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[671] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [671]),
        .Q(\f_permutation_l_/out_reg_n_0_[671] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[672] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [672]),
        .Q(\f_permutation_l_/out_reg_n_0_[672] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[673] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [673]),
        .Q(\f_permutation_l_/out_reg_n_0_[673] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[674] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [674]),
        .Q(\f_permutation_l_/out_reg_n_0_[674] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[675] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [675]),
        .Q(\f_permutation_l_/out_reg_n_0_[675] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[676] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [676]),
        .Q(\f_permutation_l_/out_reg_n_0_[676] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[677] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [677]),
        .Q(\f_permutation_l_/out_reg_n_0_[677] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[678] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [678]),
        .Q(\f_permutation_l_/out_reg_n_0_[678] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[679] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [679]),
        .Q(\f_permutation_l_/out_reg_n_0_[679] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[67] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [67]),
        .Q(\f_permutation_l_/out_reg_n_0_[67] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[680] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [680]),
        .Q(\f_permutation_l_/out_reg_n_0_[680] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[681] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [681]),
        .Q(\f_permutation_l_/out_reg_n_0_[681] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[682] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [682]),
        .Q(\f_permutation_l_/out_reg_n_0_[682] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[683] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [683]),
        .Q(\f_permutation_l_/out_reg_n_0_[683] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[684] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [684]),
        .Q(\f_permutation_l_/out_reg_n_0_[684] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[685] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [685]),
        .Q(\f_permutation_l_/out_reg_n_0_[685] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[686] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [686]),
        .Q(\f_permutation_l_/out_reg_n_0_[686] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[687] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [687]),
        .Q(\f_permutation_l_/out_reg_n_0_[687] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[688] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [688]),
        .Q(\f_permutation_l_/out_reg_n_0_[688] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[689] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [689]),
        .Q(\f_permutation_l_/out_reg_n_0_[689] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[68] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [68]),
        .Q(\f_permutation_l_/out_reg_n_0_[68] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[690] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [690]),
        .Q(\f_permutation_l_/out_reg_n_0_[690] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[691] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [691]),
        .Q(\f_permutation_l_/out_reg_n_0_[691] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[692] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [692]),
        .Q(\f_permutation_l_/out_reg_n_0_[692] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[693] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [693]),
        .Q(\f_permutation_l_/out_reg_n_0_[693] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[694] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [694]),
        .Q(\f_permutation_l_/out_reg_n_0_[694] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[695] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [695]),
        .Q(\f_permutation_l_/out_reg_n_0_[695] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[696] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [696]),
        .Q(\f_permutation_l_/out_reg_n_0_[696] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[697] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [697]),
        .Q(\f_permutation_l_/out_reg_n_0_[697] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[698] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [698]),
        .Q(\f_permutation_l_/out_reg_n_0_[698] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[699] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [699]),
        .Q(\f_permutation_l_/out_reg_n_0_[699] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[69] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [69]),
        .Q(\f_permutation_l_/out_reg_n_0_[69] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[6] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [6]),
        .Q(\f_permutation_l_/out_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[700] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [700]),
        .Q(\f_permutation_l_/out_reg_n_0_[700] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[701] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [701]),
        .Q(\f_permutation_l_/out_reg_n_0_[701] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[702] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [702]),
        .Q(\f_permutation_l_/out_reg_n_0_[702] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[703] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [703]),
        .Q(\f_permutation_l_/out_reg_n_0_[703] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[704] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [704]),
        .Q(\f_permutation_l_/out_reg_n_0_[704] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[705] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [705]),
        .Q(\f_permutation_l_/out_reg_n_0_[705] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[706] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [706]),
        .Q(\f_permutation_l_/out_reg_n_0_[706] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[707] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [707]),
        .Q(\f_permutation_l_/out_reg_n_0_[707] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[708] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [708]),
        .Q(\f_permutation_l_/out_reg_n_0_[708] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[709] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [709]),
        .Q(\f_permutation_l_/out_reg_n_0_[709] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[70] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [70]),
        .Q(\f_permutation_l_/out_reg_n_0_[70] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[710] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [710]),
        .Q(\f_permutation_l_/out_reg_n_0_[710] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[711] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [711]),
        .Q(\f_permutation_l_/out_reg_n_0_[711] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[712] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [712]),
        .Q(\f_permutation_l_/out_reg_n_0_[712] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[713] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [713]),
        .Q(\f_permutation_l_/out_reg_n_0_[713] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[714] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [714]),
        .Q(\f_permutation_l_/out_reg_n_0_[714] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[715] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [715]),
        .Q(\f_permutation_l_/out_reg_n_0_[715] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[716] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [716]),
        .Q(\f_permutation_l_/out_reg_n_0_[716] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[717] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [717]),
        .Q(\f_permutation_l_/out_reg_n_0_[717] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[718] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [718]),
        .Q(\f_permutation_l_/out_reg_n_0_[718] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[719] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [719]),
        .Q(\f_permutation_l_/out_reg_n_0_[719] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[71] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [71]),
        .Q(\f_permutation_l_/out_reg_n_0_[71] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[720] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [720]),
        .Q(\f_permutation_l_/out_reg_n_0_[720] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[721] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [721]),
        .Q(\f_permutation_l_/out_reg_n_0_[721] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[722] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [722]),
        .Q(\f_permutation_l_/out_reg_n_0_[722] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[723] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [723]),
        .Q(\f_permutation_l_/out_reg_n_0_[723] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[724] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [724]),
        .Q(\f_permutation_l_/out_reg_n_0_[724] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[725] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [725]),
        .Q(\f_permutation_l_/out_reg_n_0_[725] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[726] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [726]),
        .Q(\f_permutation_l_/out_reg_n_0_[726] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[727] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [727]),
        .Q(\f_permutation_l_/out_reg_n_0_[727] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[728] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [728]),
        .Q(\f_permutation_l_/out_reg_n_0_[728] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[729] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [729]),
        .Q(\f_permutation_l_/out_reg_n_0_[729] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[72] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [72]),
        .Q(\f_permutation_l_/out_reg_n_0_[72] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[730] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [730]),
        .Q(\f_permutation_l_/out_reg_n_0_[730] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[731] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [731]),
        .Q(\f_permutation_l_/out_reg_n_0_[731] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[732] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [732]),
        .Q(\f_permutation_l_/out_reg_n_0_[732] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[733] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [733]),
        .Q(\f_permutation_l_/out_reg_n_0_[733] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[734] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [734]),
        .Q(\f_permutation_l_/out_reg_n_0_[734] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[735] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [735]),
        .Q(\f_permutation_l_/out_reg_n_0_[735] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[736] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [736]),
        .Q(\f_permutation_l_/out_reg_n_0_[736] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[737] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [737]),
        .Q(\f_permutation_l_/out_reg_n_0_[737] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[738] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [738]),
        .Q(\f_permutation_l_/out_reg_n_0_[738] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[739] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [739]),
        .Q(\f_permutation_l_/out_reg_n_0_[739] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[73] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [73]),
        .Q(\f_permutation_l_/out_reg_n_0_[73] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[740] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [740]),
        .Q(\f_permutation_l_/out_reg_n_0_[740] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[741] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [741]),
        .Q(\f_permutation_l_/out_reg_n_0_[741] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[742] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [742]),
        .Q(\f_permutation_l_/out_reg_n_0_[742] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[743] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [743]),
        .Q(\f_permutation_l_/out_reg_n_0_[743] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[744] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [744]),
        .Q(\f_permutation_l_/out_reg_n_0_[744] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[745] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [745]),
        .Q(\f_permutation_l_/out_reg_n_0_[745] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[746] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [746]),
        .Q(\f_permutation_l_/out_reg_n_0_[746] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[747] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [747]),
        .Q(\f_permutation_l_/out_reg_n_0_[747] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[748] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [748]),
        .Q(\f_permutation_l_/out_reg_n_0_[748] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[749] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [749]),
        .Q(\f_permutation_l_/out_reg_n_0_[749] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[74] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [74]),
        .Q(\f_permutation_l_/out_reg_n_0_[74] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[750] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [750]),
        .Q(\f_permutation_l_/out_reg_n_0_[750] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[751] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [751]),
        .Q(\f_permutation_l_/out_reg_n_0_[751] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[752] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [752]),
        .Q(\f_permutation_l_/out_reg_n_0_[752] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[753] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [753]),
        .Q(\f_permutation_l_/out_reg_n_0_[753] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[754] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [754]),
        .Q(\f_permutation_l_/out_reg_n_0_[754] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[755] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [755]),
        .Q(\f_permutation_l_/out_reg_n_0_[755] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[756] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [756]),
        .Q(\f_permutation_l_/out_reg_n_0_[756] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[757] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [757]),
        .Q(\f_permutation_l_/out_reg_n_0_[757] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[758] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [758]),
        .Q(\f_permutation_l_/out_reg_n_0_[758] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[759] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [759]),
        .Q(\f_permutation_l_/out_reg_n_0_[759] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[75] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [75]),
        .Q(\f_permutation_l_/out_reg_n_0_[75] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[760] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [760]),
        .Q(\f_permutation_l_/out_reg_n_0_[760] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[761] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [761]),
        .Q(\f_permutation_l_/out_reg_n_0_[761] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[762] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [762]),
        .Q(\f_permutation_l_/out_reg_n_0_[762] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[763] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [763]),
        .Q(\f_permutation_l_/out_reg_n_0_[763] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[764] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [764]),
        .Q(\f_permutation_l_/out_reg_n_0_[764] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[765] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [765]),
        .Q(\f_permutation_l_/out_reg_n_0_[765] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[766] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [766]),
        .Q(\f_permutation_l_/out_reg_n_0_[766] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[767] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [767]),
        .Q(\f_permutation_l_/out_reg_n_0_[767] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[768] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [768]),
        .Q(\f_permutation_l_/out_reg_n_0_[768] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[769] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [769]),
        .Q(\f_permutation_l_/out_reg_n_0_[769] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[76] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [76]),
        .Q(\f_permutation_l_/out_reg_n_0_[76] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[770] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [770]),
        .Q(\f_permutation_l_/out_reg_n_0_[770] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[771] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [771]),
        .Q(\f_permutation_l_/out_reg_n_0_[771] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[772] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [772]),
        .Q(\f_permutation_l_/out_reg_n_0_[772] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[773] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [773]),
        .Q(\f_permutation_l_/out_reg_n_0_[773] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[774] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [774]),
        .Q(\f_permutation_l_/out_reg_n_0_[774] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[775] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [775]),
        .Q(\f_permutation_l_/out_reg_n_0_[775] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[776] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [776]),
        .Q(\f_permutation_l_/out_reg_n_0_[776] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[777] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [777]),
        .Q(\f_permutation_l_/out_reg_n_0_[777] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[778] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [778]),
        .Q(\f_permutation_l_/out_reg_n_0_[778] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[779] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [779]),
        .Q(\f_permutation_l_/out_reg_n_0_[779] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[77] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [77]),
        .Q(\f_permutation_l_/out_reg_n_0_[77] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[780] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [780]),
        .Q(\f_permutation_l_/out_reg_n_0_[780] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[781] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [781]),
        .Q(\f_permutation_l_/out_reg_n_0_[781] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[782] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [782]),
        .Q(\f_permutation_l_/out_reg_n_0_[782] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[783] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [783]),
        .Q(\f_permutation_l_/out_reg_n_0_[783] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[784] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [784]),
        .Q(\f_permutation_l_/out_reg_n_0_[784] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[785] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [785]),
        .Q(\f_permutation_l_/out_reg_n_0_[785] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[786] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [786]),
        .Q(\f_permutation_l_/out_reg_n_0_[786] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[787] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [787]),
        .Q(\f_permutation_l_/out_reg_n_0_[787] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[788] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [788]),
        .Q(\f_permutation_l_/out_reg_n_0_[788] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[789] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [789]),
        .Q(\f_permutation_l_/out_reg_n_0_[789] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[78] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [78]),
        .Q(\f_permutation_l_/out_reg_n_0_[78] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[790] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [790]),
        .Q(\f_permutation_l_/out_reg_n_0_[790] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[791] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [791]),
        .Q(\f_permutation_l_/out_reg_n_0_[791] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[792] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [792]),
        .Q(\f_permutation_l_/out_reg_n_0_[792] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[793] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [793]),
        .Q(\f_permutation_l_/out_reg_n_0_[793] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[794] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [794]),
        .Q(\f_permutation_l_/out_reg_n_0_[794] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[795] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [795]),
        .Q(\f_permutation_l_/out_reg_n_0_[795] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[796] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [796]),
        .Q(\f_permutation_l_/out_reg_n_0_[796] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[797] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [797]),
        .Q(\f_permutation_l_/out_reg_n_0_[797] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[798] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [798]),
        .Q(\f_permutation_l_/out_reg_n_0_[798] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[799] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [799]),
        .Q(\f_permutation_l_/out_reg_n_0_[799] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[79] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [79]),
        .Q(\f_permutation_l_/out_reg_n_0_[79] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[7] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [7]),
        .Q(\f_permutation_l_/out_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[800] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [800]),
        .Q(\f_permutation_l_/out_reg_n_0_[800] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[801] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [801]),
        .Q(\f_permutation_l_/out_reg_n_0_[801] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[802] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [802]),
        .Q(\f_permutation_l_/out_reg_n_0_[802] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[803] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [803]),
        .Q(\f_permutation_l_/out_reg_n_0_[803] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[804] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [804]),
        .Q(\f_permutation_l_/out_reg_n_0_[804] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[805] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [805]),
        .Q(\f_permutation_l_/out_reg_n_0_[805] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[806] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [806]),
        .Q(\f_permutation_l_/out_reg_n_0_[806] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[807] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [807]),
        .Q(\f_permutation_l_/out_reg_n_0_[807] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[808] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [808]),
        .Q(\f_permutation_l_/out_reg_n_0_[808] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[809] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [809]),
        .Q(\f_permutation_l_/out_reg_n_0_[809] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[80] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [80]),
        .Q(\f_permutation_l_/out_reg_n_0_[80] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[810] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [810]),
        .Q(\f_permutation_l_/out_reg_n_0_[810] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[811] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [811]),
        .Q(\f_permutation_l_/out_reg_n_0_[811] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[812] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [812]),
        .Q(\f_permutation_l_/out_reg_n_0_[812] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[813] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [813]),
        .Q(\f_permutation_l_/out_reg_n_0_[813] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[814] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [814]),
        .Q(\f_permutation_l_/out_reg_n_0_[814] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[815] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [815]),
        .Q(\f_permutation_l_/out_reg_n_0_[815] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[816] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [816]),
        .Q(\f_permutation_l_/out_reg_n_0_[816] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[817] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [817]),
        .Q(\f_permutation_l_/out_reg_n_0_[817] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[818] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [818]),
        .Q(\f_permutation_l_/out_reg_n_0_[818] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[819] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [819]),
        .Q(\f_permutation_l_/out_reg_n_0_[819] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[81] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [81]),
        .Q(\f_permutation_l_/out_reg_n_0_[81] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[820] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [820]),
        .Q(\f_permutation_l_/out_reg_n_0_[820] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[821] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [821]),
        .Q(\f_permutation_l_/out_reg_n_0_[821] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[822] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [822]),
        .Q(\f_permutation_l_/out_reg_n_0_[822] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[823] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [823]),
        .Q(\f_permutation_l_/out_reg_n_0_[823] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[824] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [824]),
        .Q(\f_permutation_l_/out_reg_n_0_[824] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[825] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [825]),
        .Q(\f_permutation_l_/out_reg_n_0_[825] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[826] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [826]),
        .Q(\f_permutation_l_/out_reg_n_0_[826] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[827] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [827]),
        .Q(\f_permutation_l_/out_reg_n_0_[827] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[828] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [828]),
        .Q(\f_permutation_l_/out_reg_n_0_[828] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[829] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [829]),
        .Q(\f_permutation_l_/out_reg_n_0_[829] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[82] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [82]),
        .Q(\f_permutation_l_/out_reg_n_0_[82] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[830] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [830]),
        .Q(\f_permutation_l_/out_reg_n_0_[830] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[831] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [831]),
        .Q(\f_permutation_l_/out_reg_n_0_[831] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[832] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [832]),
        .Q(\f_permutation_l_/out_reg_n_0_[832] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[833] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [833]),
        .Q(\f_permutation_l_/out_reg_n_0_[833] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[834] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [834]),
        .Q(\f_permutation_l_/out_reg_n_0_[834] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[835] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [835]),
        .Q(\f_permutation_l_/out_reg_n_0_[835] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[836] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [836]),
        .Q(\f_permutation_l_/out_reg_n_0_[836] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[837] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [837]),
        .Q(\f_permutation_l_/out_reg_n_0_[837] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[838] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [838]),
        .Q(\f_permutation_l_/out_reg_n_0_[838] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[839] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [839]),
        .Q(\f_permutation_l_/out_reg_n_0_[839] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[83] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [83]),
        .Q(\f_permutation_l_/out_reg_n_0_[83] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[840] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [840]),
        .Q(\f_permutation_l_/out_reg_n_0_[840] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[841] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [841]),
        .Q(\f_permutation_l_/out_reg_n_0_[841] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[842] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [842]),
        .Q(\f_permutation_l_/out_reg_n_0_[842] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[843] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [843]),
        .Q(\f_permutation_l_/out_reg_n_0_[843] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[844] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [844]),
        .Q(\f_permutation_l_/out_reg_n_0_[844] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[845] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [845]),
        .Q(\f_permutation_l_/out_reg_n_0_[845] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[846] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [846]),
        .Q(\f_permutation_l_/out_reg_n_0_[846] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[847] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [847]),
        .Q(\f_permutation_l_/out_reg_n_0_[847] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[848] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [848]),
        .Q(\f_permutation_l_/out_reg_n_0_[848] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[849] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [849]),
        .Q(\f_permutation_l_/out_reg_n_0_[849] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[84] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [84]),
        .Q(\f_permutation_l_/out_reg_n_0_[84] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[850] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [850]),
        .Q(\f_permutation_l_/out_reg_n_0_[850] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[851] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [851]),
        .Q(\f_permutation_l_/out_reg_n_0_[851] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[852] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [852]),
        .Q(\f_permutation_l_/out_reg_n_0_[852] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[853] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [853]),
        .Q(\f_permutation_l_/out_reg_n_0_[853] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[854] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [854]),
        .Q(\f_permutation_l_/out_reg_n_0_[854] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[855] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [855]),
        .Q(\f_permutation_l_/out_reg_n_0_[855] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[856] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [856]),
        .Q(\f_permutation_l_/out_reg_n_0_[856] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[857] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [857]),
        .Q(\f_permutation_l_/out_reg_n_0_[857] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[858] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [858]),
        .Q(\f_permutation_l_/out_reg_n_0_[858] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[859] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [859]),
        .Q(\f_permutation_l_/out_reg_n_0_[859] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[85] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [85]),
        .Q(\f_permutation_l_/out_reg_n_0_[85] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[860] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [860]),
        .Q(\f_permutation_l_/out_reg_n_0_[860] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[861] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [861]),
        .Q(\f_permutation_l_/out_reg_n_0_[861] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[862] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [862]),
        .Q(\f_permutation_l_/out_reg_n_0_[862] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[863] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [863]),
        .Q(\f_permutation_l_/out_reg_n_0_[863] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[864] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [864]),
        .Q(\f_permutation_l_/out_reg_n_0_[864] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[865] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [865]),
        .Q(\f_permutation_l_/out_reg_n_0_[865] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[866] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [866]),
        .Q(\f_permutation_l_/out_reg_n_0_[866] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[867] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [867]),
        .Q(\f_permutation_l_/out_reg_n_0_[867] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[868] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [868]),
        .Q(\f_permutation_l_/out_reg_n_0_[868] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[869] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [869]),
        .Q(\f_permutation_l_/out_reg_n_0_[869] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[86] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [86]),
        .Q(\f_permutation_l_/out_reg_n_0_[86] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[870] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [870]),
        .Q(\f_permutation_l_/out_reg_n_0_[870] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[871] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [871]),
        .Q(\f_permutation_l_/out_reg_n_0_[871] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[872] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [872]),
        .Q(\f_permutation_l_/out_reg_n_0_[872] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[873] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [873]),
        .Q(\f_permutation_l_/out_reg_n_0_[873] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[874] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [874]),
        .Q(\f_permutation_l_/out_reg_n_0_[874] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[875] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [875]),
        .Q(\f_permutation_l_/out_reg_n_0_[875] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[876] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [876]),
        .Q(\f_permutation_l_/out_reg_n_0_[876] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[877] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [877]),
        .Q(\f_permutation_l_/out_reg_n_0_[877] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[878] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [878]),
        .Q(\f_permutation_l_/out_reg_n_0_[878] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[879] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [879]),
        .Q(\f_permutation_l_/out_reg_n_0_[879] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[87] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [87]),
        .Q(\f_permutation_l_/out_reg_n_0_[87] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[880] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [880]),
        .Q(\f_permutation_l_/out_reg_n_0_[880] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[881] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [881]),
        .Q(\f_permutation_l_/out_reg_n_0_[881] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[882] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [882]),
        .Q(\f_permutation_l_/out_reg_n_0_[882] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[883] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [883]),
        .Q(\f_permutation_l_/out_reg_n_0_[883] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[884] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [884]),
        .Q(\f_permutation_l_/out_reg_n_0_[884] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[885] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [885]),
        .Q(\f_permutation_l_/out_reg_n_0_[885] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[886] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [886]),
        .Q(\f_permutation_l_/out_reg_n_0_[886] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[887] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [887]),
        .Q(\f_permutation_l_/out_reg_n_0_[887] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[888] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [888]),
        .Q(\f_permutation_l_/out_reg_n_0_[888] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[889] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [889]),
        .Q(\f_permutation_l_/out_reg_n_0_[889] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[88] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [88]),
        .Q(\f_permutation_l_/out_reg_n_0_[88] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[890] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [890]),
        .Q(\f_permutation_l_/out_reg_n_0_[890] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[891] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [891]),
        .Q(\f_permutation_l_/out_reg_n_0_[891] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[892] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [892]),
        .Q(\f_permutation_l_/out_reg_n_0_[892] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[893] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [893]),
        .Q(\f_permutation_l_/out_reg_n_0_[893] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[894] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [894]),
        .Q(\f_permutation_l_/out_reg_n_0_[894] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[895] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [895]),
        .Q(\f_permutation_l_/out_reg_n_0_[895] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[896] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [896]),
        .Q(\f_permutation_l_/out_reg_n_0_[896] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[897] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [897]),
        .Q(\f_permutation_l_/out_reg_n_0_[897] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[898] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [898]),
        .Q(\f_permutation_l_/out_reg_n_0_[898] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[899] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [899]),
        .Q(\f_permutation_l_/out_reg_n_0_[899] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[89] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [89]),
        .Q(\f_permutation_l_/out_reg_n_0_[89] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[8] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [8]),
        .Q(\f_permutation_l_/out_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[900] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [900]),
        .Q(\f_permutation_l_/out_reg_n_0_[900] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[901] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [901]),
        .Q(\f_permutation_l_/out_reg_n_0_[901] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[902] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [902]),
        .Q(\f_permutation_l_/out_reg_n_0_[902] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[903] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [903]),
        .Q(\f_permutation_l_/out_reg_n_0_[903] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[904] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [904]),
        .Q(\f_permutation_l_/out_reg_n_0_[904] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[905] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [905]),
        .Q(\f_permutation_l_/out_reg_n_0_[905] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[906] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [906]),
        .Q(\f_permutation_l_/out_reg_n_0_[906] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[907] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [907]),
        .Q(\f_permutation_l_/out_reg_n_0_[907] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[908] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [908]),
        .Q(\f_permutation_l_/out_reg_n_0_[908] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[909] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [909]),
        .Q(\f_permutation_l_/out_reg_n_0_[909] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[90] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [90]),
        .Q(\f_permutation_l_/out_reg_n_0_[90] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[910] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [910]),
        .Q(\f_permutation_l_/out_reg_n_0_[910] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[911] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [911]),
        .Q(\f_permutation_l_/out_reg_n_0_[911] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[912] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [912]),
        .Q(\f_permutation_l_/out_reg_n_0_[912] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[913] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [913]),
        .Q(\f_permutation_l_/out_reg_n_0_[913] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[914] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [914]),
        .Q(\f_permutation_l_/out_reg_n_0_[914] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[915] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [915]),
        .Q(\f_permutation_l_/out_reg_n_0_[915] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[916] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [916]),
        .Q(\f_permutation_l_/out_reg_n_0_[916] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[917] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [917]),
        .Q(\f_permutation_l_/out_reg_n_0_[917] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[918] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [918]),
        .Q(\f_permutation_l_/out_reg_n_0_[918] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[919] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [919]),
        .Q(\f_permutation_l_/out_reg_n_0_[919] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[91] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [91]),
        .Q(\f_permutation_l_/out_reg_n_0_[91] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[920] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [920]),
        .Q(\f_permutation_l_/out_reg_n_0_[920] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[921] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [921]),
        .Q(\f_permutation_l_/out_reg_n_0_[921] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[922] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [922]),
        .Q(\f_permutation_l_/out_reg_n_0_[922] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[923] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [923]),
        .Q(\f_permutation_l_/out_reg_n_0_[923] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[924] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [924]),
        .Q(\f_permutation_l_/out_reg_n_0_[924] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[925] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [925]),
        .Q(\f_permutation_l_/out_reg_n_0_[925] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[926] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [926]),
        .Q(\f_permutation_l_/out_reg_n_0_[926] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[927] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [927]),
        .Q(\f_permutation_l_/out_reg_n_0_[927] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[928] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [928]),
        .Q(\f_permutation_l_/out_reg_n_0_[928] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[929] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [929]),
        .Q(\f_permutation_l_/out_reg_n_0_[929] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[92] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [92]),
        .Q(\f_permutation_l_/out_reg_n_0_[92] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[930] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [930]),
        .Q(\f_permutation_l_/out_reg_n_0_[930] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[931] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [931]),
        .Q(\f_permutation_l_/out_reg_n_0_[931] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[932] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [932]),
        .Q(\f_permutation_l_/out_reg_n_0_[932] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[933] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [933]),
        .Q(\f_permutation_l_/out_reg_n_0_[933] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[934] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [934]),
        .Q(\f_permutation_l_/out_reg_n_0_[934] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[935] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [935]),
        .Q(\f_permutation_l_/out_reg_n_0_[935] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[936] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [936]),
        .Q(\f_permutation_l_/out_reg_n_0_[936] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[937] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [937]),
        .Q(\f_permutation_l_/out_reg_n_0_[937] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[938] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [938]),
        .Q(\f_permutation_l_/out_reg_n_0_[938] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[939] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [939]),
        .Q(\f_permutation_l_/out_reg_n_0_[939] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[93] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [93]),
        .Q(\f_permutation_l_/out_reg_n_0_[93] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[940] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [940]),
        .Q(\f_permutation_l_/out_reg_n_0_[940] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[941] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [941]),
        .Q(\f_permutation_l_/out_reg_n_0_[941] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[942] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [942]),
        .Q(\f_permutation_l_/out_reg_n_0_[942] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[943] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [943]),
        .Q(\f_permutation_l_/out_reg_n_0_[943] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[944] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [944]),
        .Q(\f_permutation_l_/out_reg_n_0_[944] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[945] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [945]),
        .Q(\f_permutation_l_/out_reg_n_0_[945] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[946] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [946]),
        .Q(\f_permutation_l_/out_reg_n_0_[946] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[947] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [947]),
        .Q(\f_permutation_l_/out_reg_n_0_[947] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[948] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [948]),
        .Q(\f_permutation_l_/out_reg_n_0_[948] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[949] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [949]),
        .Q(\f_permutation_l_/out_reg_n_0_[949] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[94] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [94]),
        .Q(\f_permutation_l_/out_reg_n_0_[94] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[950] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [950]),
        .Q(\f_permutation_l_/out_reg_n_0_[950] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[951] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [951]),
        .Q(\f_permutation_l_/out_reg_n_0_[951] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[952] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [952]),
        .Q(\f_permutation_l_/out_reg_n_0_[952] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[953] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [953]),
        .Q(\f_permutation_l_/out_reg_n_0_[953] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[954] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [954]),
        .Q(\f_permutation_l_/out_reg_n_0_[954] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[955] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [955]),
        .Q(\f_permutation_l_/out_reg_n_0_[955] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[956] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [956]),
        .Q(\f_permutation_l_/out_reg_n_0_[956] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[957] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [957]),
        .Q(\f_permutation_l_/out_reg_n_0_[957] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[958] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [958]),
        .Q(\f_permutation_l_/out_reg_n_0_[958] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[959] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [959]),
        .Q(\f_permutation_l_/out_reg_n_0_[959] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[95] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [95]),
        .Q(\f_permutation_l_/out_reg_n_0_[95] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[960] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [960]),
        .Q(\f_permutation_l_/out_reg_n_0_[960] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[961] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [961]),
        .Q(\f_permutation_l_/out_reg_n_0_[961] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[962] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [962]),
        .Q(\f_permutation_l_/out_reg_n_0_[962] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[963] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [963]),
        .Q(\f_permutation_l_/out_reg_n_0_[963] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[964] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [964]),
        .Q(\f_permutation_l_/out_reg_n_0_[964] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[965] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [965]),
        .Q(\f_permutation_l_/out_reg_n_0_[965] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[966] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [966]),
        .Q(\f_permutation_l_/out_reg_n_0_[966] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[967] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [967]),
        .Q(\f_permutation_l_/out_reg_n_0_[967] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[968] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [968]),
        .Q(\f_permutation_l_/out_reg_n_0_[968] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[969] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [969]),
        .Q(\f_permutation_l_/out_reg_n_0_[969] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[96] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [96]),
        .Q(\f_permutation_l_/out_reg_n_0_[96] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[970] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [970]),
        .Q(\f_permutation_l_/out_reg_n_0_[970] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[971] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [971]),
        .Q(\f_permutation_l_/out_reg_n_0_[971] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[972] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [972]),
        .Q(\f_permutation_l_/out_reg_n_0_[972] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[973] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [973]),
        .Q(\f_permutation_l_/out_reg_n_0_[973] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[974] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [974]),
        .Q(\f_permutation_l_/out_reg_n_0_[974] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[975] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [975]),
        .Q(\f_permutation_l_/out_reg_n_0_[975] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[976] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [976]),
        .Q(\f_permutation_l_/out_reg_n_0_[976] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[977] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [977]),
        .Q(\f_permutation_l_/out_reg_n_0_[977] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[978] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [978]),
        .Q(\f_permutation_l_/out_reg_n_0_[978] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[979] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [979]),
        .Q(\f_permutation_l_/out_reg_n_0_[979] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[97] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [97]),
        .Q(\f_permutation_l_/out_reg_n_0_[97] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[980] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [980]),
        .Q(\f_permutation_l_/out_reg_n_0_[980] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[981] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [981]),
        .Q(\f_permutation_l_/out_reg_n_0_[981] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[982] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [982]),
        .Q(\f_permutation_l_/out_reg_n_0_[982] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[983] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [983]),
        .Q(\f_permutation_l_/out_reg_n_0_[983] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[984] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [984]),
        .Q(\f_permutation_l_/out_reg_n_0_[984] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[985] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [985]),
        .Q(\f_permutation_l_/out_reg_n_0_[985] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[986] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [986]),
        .Q(\f_permutation_l_/out_reg_n_0_[986] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[987] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [987]),
        .Q(\f_permutation_l_/out_reg_n_0_[987] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[988] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [988]),
        .Q(\f_permutation_l_/out_reg_n_0_[988] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[989] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [989]),
        .Q(\f_permutation_l_/out_reg_n_0_[989] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[98] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [98]),
        .Q(\f_permutation_l_/out_reg_n_0_[98] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[990] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [990]),
        .Q(\f_permutation_l_/out_reg_n_0_[990] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[991] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [991]),
        .Q(\f_permutation_l_/out_reg_n_0_[991] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[992] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [992]),
        .Q(\f_permutation_l_/out_reg_n_0_[992] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[993] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [993]),
        .Q(\f_permutation_l_/out_reg_n_0_[993] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[994] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [994]),
        .Q(\f_permutation_l_/out_reg_n_0_[994] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[995] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [995]),
        .Q(\f_permutation_l_/out_reg_n_0_[995] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[996] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [996]),
        .Q(\f_permutation_l_/out_reg_n_0_[996] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[997] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [997]),
        .Q(\f_permutation_l_/out_reg_n_0_[997] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[998] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [998]),
        .Q(\f_permutation_l_/out_reg_n_0_[998] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[999] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [999]),
        .Q(\f_permutation_l_/out_reg_n_0_[999] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[99] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [99]),
        .Q(\f_permutation_l_/out_reg_n_0_[99] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \f_permutation_l_/out_reg[9] 
       (.C(clk),
        .CE(\f_permutation_l_/update ),
        .D(\f_permutation_l_/round_out [9]),
        .Q(\f_permutation_l_/out_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \i[0]_i_1 
       (.I0(\f_permutation_l_/calc ),
        .I1(buffer_full),
        .O(\i[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[0]_i_1__0 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\i[0]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[10]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[9] ),
        .I1(update__0_i_1_n_0),
        .O(\i[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[11]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[10] ),
        .I1(update__0_i_1_n_0),
        .O(\i[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[12]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[11] ),
        .I1(update__0_i_1_n_0),
        .O(\i[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[13]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[12] ),
        .I1(update__0_i_1_n_0),
        .O(\i[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[14]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[13] ),
        .I1(update__0_i_1_n_0),
        .O(\i[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[15]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[14] ),
        .I1(update__0_i_1_n_0),
        .O(\i[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[16]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[15] ),
        .I1(update__0_i_1_n_0),
        .O(\i[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[17]_i_1 
       (.I0(\padder_l_/p_0_in ),
        .I1(update__0_i_1_n_0),
        .O(\i[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair302" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[1]_i_1 
       (.I0(\padder_l_/i_reg_n_0_ ),
        .I1(update__0_i_1_n_0),
        .O(\i[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair303" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[2]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[1] ),
        .I1(update__0_i_1_n_0),
        .O(\i[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair304" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[3]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[2] ),
        .I1(update__0_i_1_n_0),
        .O(\i[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair305" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[4]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[3] ),
        .I1(update__0_i_1_n_0),
        .O(\i[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair306" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[5]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[4] ),
        .I1(update__0_i_1_n_0),
        .O(\i[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair307" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[6]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[5] ),
        .I1(update__0_i_1_n_0),
        .O(\i[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair308" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[7]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[6] ),
        .I1(update__0_i_1_n_0),
        .O(\i[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair309" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[8]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[7] ),
        .I1(update__0_i_1_n_0),
        .O(\i[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \i[9]_i_1 
       (.I0(\padder_l_/i_reg_n_0_[8] ),
        .I1(update__0_i_1_n_0),
        .O(\i[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "sha3_low_throughput_0/\i_reg " *) 
  (* srl_name = "sha3_low_throughput_0/\i_reg[20]_srl21___i_reg_r_19 " *) 
  SRLC32E #(
    .INIT(32'h00000000),
    .IS_CLK_INVERTED(1'b0)) 
    \i_reg[20]_srl21___i_reg_r_19 
       (.A({\<const1>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(p_0_out),
        .Q(i_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \i_reg[20]_srl21___i_reg_r_19_i_1 
       (.I0(\i[0]_i_1__0_n_0 ),
        .I1(state),
        .O(p_0_out));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \i_reg[21]_i_reg_r_20 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg),
        .Q(\i_reg[21]_i_reg_r_20_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \i_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_gate_n_0),
        .Q(i),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    i_reg_gate
       (.I0(\i_reg[21]_i_reg_r_20_n_0 ),
        .I1(i_reg_r_20_n_0),
        .O(i_reg_gate_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\<const1>__0__0 ),
        .Q(i_reg_r_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_0
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_n_0),
        .Q(i_reg_r_0_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_1
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_0_n_0),
        .Q(i_reg_r_1_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_10
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_9_n_0),
        .Q(i_reg_r_10_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_11
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_10_n_0),
        .Q(i_reg_r_11_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_12
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_11_n_0),
        .Q(i_reg_r_12_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_13
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_12_n_0),
        .Q(i_reg_r_13_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_14
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_13_n_0),
        .Q(i_reg_r_14_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_15
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_14_n_0),
        .Q(i_reg_r_15_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_16
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_15_n_0),
        .Q(i_reg_r_16_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_17
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_16_n_0),
        .Q(i_reg_r_17_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_18
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_17_n_0),
        .Q(i_reg_r_18_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_19
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_18_n_0),
        .Q(i_reg_r_19_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_2
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_1_n_0),
        .Q(i_reg_r_2_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_20
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_19_n_0),
        .Q(i_reg_r_20_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_3
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_2_n_0),
        .Q(i_reg_r_3_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_4
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_3_n_0),
        .Q(i_reg_r_4_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_5
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_4_n_0),
        .Q(i_reg_r_5_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_6
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_5_n_0),
        .Q(i_reg_r_6_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_7
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_6_n_0),
        .Q(i_reg_r_7_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_8
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_7_n_0),
        .Q(i_reg_r_8_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    i_reg_r_9
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(i_reg_r_8_n_0),
        .Q(i_reg_r_9_n_0),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[0]_i_1 
       (.I0(\out[1578]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[254] ),
        .I2(\out[256]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1033]),
        .I4(\out[1502]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1000]_i_1 
       (.I0(\out[1558]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[171] ),
        .I2(\out[1256]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[980] ),
        .I4(\out[1442]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1000]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1001]_i_1 
       (.I0(\out[1559]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[172] ),
        .I2(\out[1257]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[981] ),
        .I4(\out[1443]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1001]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1002]_i_1 
       (.I0(\out[1560]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[173] ),
        .I2(\out[1258]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[982] ),
        .I4(\out[1444]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1002]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1003]_i_1 
       (.I0(\out[1561]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[174] ),
        .I2(\out[1259]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[983] ),
        .I4(\out[1445]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1003]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1004]_i_1 
       (.I0(\out[1562]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[175] ),
        .I2(\out[1260]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[984] ),
        .I4(\out[1446]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1004]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1005]_i_1 
       (.I0(\out[1563]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[176] ),
        .I2(\out[1261]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[985] ),
        .I4(\out[1447]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1005]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1006]_i_1 
       (.I0(\out[1564]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[177] ),
        .I2(\out[1262]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[986] ),
        .I4(\out[1448]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1006]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1007]_i_1 
       (.I0(\out[1565]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[178] ),
        .I2(\out[1263]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[987] ),
        .I4(\out[1449]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1007]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1008]_i_1 
       (.I0(\out[1566]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[179] ),
        .I2(\out[1264]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[988] ),
        .I4(\out[1450]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1008]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1009]_i_1 
       (.I0(\out[1567]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[180] ),
        .I2(\out[1265]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[989] ),
        .I4(\out[1451]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1009]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[100]_i_1 
       (.I0(\out[1278]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[635] ),
        .I2(\f_permutation_l_/out_reg_n_0_[226] ),
        .I3(\out[1550]_i_3_n_0 ),
        .I4(\out[292]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1010]_i_1 
       (.I0(\out[1568]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[181] ),
        .I2(\out[1266]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[990] ),
        .I4(\out[1452]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1010]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1011]_i_1 
       (.I0(\out[1569]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[182] ),
        .I2(\out[1267]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[991] ),
        .I4(\out[1453]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1011]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1012]_i_1 
       (.I0(\out[1570]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[183] ),
        .I2(\out[1268]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[992] ),
        .I4(\out[1454]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1012]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1013]_i_1 
       (.I0(\out[1571]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[184] ),
        .I2(\out[1269]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[993] ),
        .I4(\out[1455]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1013]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1014]_i_1 
       (.I0(\out[1572]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[185] ),
        .I2(\out[1270]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[994] ),
        .I4(\out[1456]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1014]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1015]_i_1 
       (.I0(\out[1573]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[186] ),
        .I2(\out[1271]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[995] ),
        .I4(\out[1457]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1015]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1016]_i_1 
       (.I0(\out[1574]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[187] ),
        .I2(\out[1272]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[996] ),
        .I4(\out[1458]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1016]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1017]_i_1 
       (.I0(\out[1575]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[188] ),
        .I2(\out[1273]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[997] ),
        .I4(\out[1459]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1017]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1018]_i_1 
       (.I0(\out[1576]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[189] ),
        .I2(\out[1274]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[998] ),
        .I4(\out[1460]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1018]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1019]_i_1 
       (.I0(\out[1577]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[190] ),
        .I2(\out[1275]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[999] ),
        .I4(\out[1461]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1019]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[101]_i_1 
       (.I0(\out[1279]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[636] ),
        .I2(\f_permutation_l_/out_reg_n_0_[227] ),
        .I3(\out[1295]_i_3_n_0 ),
        .I4(\out[293]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1020]_i_1 
       (.I0(\out[1578]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[191] ),
        .I2(\out[1276]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1000] ),
        .I4(\out[1462]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1020]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1021]_i_1 
       (.I0(\out[1579]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[128] ),
        .I2(\out[1277]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1001] ),
        .I4(\out[1463]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1021]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1022]_i_1 
       (.I0(\out[1580]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[129] ),
        .I2(\out[1278]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1002] ),
        .I4(\out[1464]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1022]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1023]_i_1 
       (.I0(\out[1581]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[130] ),
        .I2(\out[1279]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1003] ),
        .I4(\out[1465]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1023]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1024]_i_1 
       (.I0(\out[1343]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[531] ),
        .I2(\f_permutation_l_/out_reg_n_0_[131] ),
        .I3(\out[1582]_i_4_n_0 ),
        .I4(\out[1216]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1024]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1025]_i_1 
       (.I0(\out[1280]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[532] ),
        .I2(\f_permutation_l_/out_reg_n_0_[132] ),
        .I3(\out[1583]_i_4_n_0 ),
        .I4(\out[1217]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1025]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1026]_i_1 
       (.I0(\out[1281]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[533] ),
        .I2(\f_permutation_l_/out_reg_n_0_[133] ),
        .I3(\out[1584]_i_4_n_0 ),
        .I4(\out[1218]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1026]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1027]_i_1 
       (.I0(\out[1538]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[534] ),
        .I2(\f_permutation_l_/out_reg_n_0_[134] ),
        .I3(\out[1585]_i_4_n_0 ),
        .I4(\out[1219]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1027]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1028]_i_1 
       (.I0(\out[1539]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[535] ),
        .I2(\f_permutation_l_/out_reg_n_0_[135] ),
        .I3(\out[1586]_i_4_n_0 ),
        .I4(\out[1220]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1028]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1029]_i_1 
       (.I0(\out[1540]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[536] ),
        .I2(\f_permutation_l_/out_reg_n_0_[136] ),
        .I3(\out[1587]_i_4_n_0 ),
        .I4(\out[1221]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1029]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[102]_i_1 
       (.I0(\out[1216]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[637] ),
        .I2(\f_permutation_l_/out_reg_n_0_[228] ),
        .I3(\out[1552]_i_3_n_0 ),
        .I4(\out[294]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1030]_i_1 
       (.I0(\out[1541]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[537] ),
        .I2(\f_permutation_l_/out_reg_n_0_[137] ),
        .I3(\out[1588]_i_4_n_0 ),
        .I4(\out[1222]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1030]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1031]_i_1 
       (.I0(\out[1542]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[538] ),
        .I2(\f_permutation_l_/out_reg_n_0_[138] ),
        .I3(\out[1589]_i_4_n_0 ),
        .I4(\out[1223]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1031]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1032]_i_1 
       (.I0(\out[1287]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[539] ),
        .I2(\f_permutation_l_/out_reg_n_0_[139] ),
        .I3(\out[1590]_i_4_n_0 ),
        .I4(\out[1224]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1032]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1033]_i_1 
       (.I0(\out[1544]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[540] ),
        .I2(\f_permutation_l_/out_reg_n_0_[140] ),
        .I3(\out[1591]_i_4_n_0 ),
        .I4(\out[1225]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1033]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1034]_i_1 
       (.I0(\out[1545]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[541] ),
        .I2(\f_permutation_l_/out_reg_n_0_[141] ),
        .I3(\out[1592]_i_4_n_0 ),
        .I4(\out[1226]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1034]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1035]_i_1 
       (.I0(\out[1546]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[542] ),
        .I2(\f_permutation_l_/out_reg_n_0_[142] ),
        .I3(\out[1593]_i_4_n_0 ),
        .I4(\out[1227]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1035]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1036]_i_1 
       (.I0(\out[1547]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[543] ),
        .I2(\f_permutation_l_/out_reg_n_0_[143] ),
        .I3(\out[1594]_i_4_n_0 ),
        .I4(\out[1228]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1036]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1037]_i_1 
       (.I0(\out[1548]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[544] ),
        .I2(\f_permutation_l_/out_reg_n_0_[144] ),
        .I3(\out[1595]_i_4_n_0 ),
        .I4(\out[1229]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1037]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1038]_i_1 
       (.I0(\out[1549]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[545] ),
        .I2(\f_permutation_l_/out_reg_n_0_[145] ),
        .I3(\out[1596]_i_4_n_0 ),
        .I4(\out[1230]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1038]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1039]_i_1 
       (.I0(\out[1550]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[546] ),
        .I2(\f_permutation_l_/out_reg_n_0_[146] ),
        .I3(\out[1597]_i_4_n_0 ),
        .I4(\out[1231]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1039]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[103]_i_1 
       (.I0(\out[1217]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[638] ),
        .I2(\f_permutation_l_/out_reg_n_0_[229] ),
        .I3(\out[1553]_i_3_n_0 ),
        .I4(\out[295]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1040]_i_1 
       (.I0(\out[1295]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[547] ),
        .I2(\f_permutation_l_/out_reg_n_0_[147] ),
        .I3(\out[1598]_i_4_n_0 ),
        .I4(\out[1232]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1040]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1041]_i_1 
       (.I0(\out[1552]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[548] ),
        .I2(\f_permutation_l_/out_reg_n_0_[148] ),
        .I3(\out[1599]_i_3_n_0 ),
        .I4(\out[1233]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1041]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1042]_i_1 
       (.I0(\out[1553]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[549] ),
        .I2(\f_permutation_l_/out_reg_n_0_[149] ),
        .I3(\out[1472]_i_2_n_0 ),
        .I4(\out[1234]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1042]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1043]_i_1 
       (.I0(\out[1554]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[550] ),
        .I2(\f_permutation_l_/out_reg_n_0_[150] ),
        .I3(\out[1537]_i_3_n_0 ),
        .I4(\out[1235]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1043]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1044]_i_1 
       (.I0(\out[1555]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[551] ),
        .I2(\f_permutation_l_/out_reg_n_0_[151] ),
        .I3(\out[1538]_i_4_n_0 ),
        .I4(\out[1236]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1044]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1045]_i_1 
       (.I0(\out[1556]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[552] ),
        .I2(\f_permutation_l_/out_reg_n_0_[152] ),
        .I3(\out[1045]_i_2_n_0 ),
        .I4(\out[1237]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1045]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1045]_i_2 
       (.I0(\out[1539]_i_14_n_0 ),
        .I1(padder_out_1[480]),
        .I2(out[416]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\f_permutation_l_/round_in [1367]),
        .I5(\out[1539]_i_12_n_0 ),
        .O(\out[1045]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1046]_i_1 
       (.I0(\out[1557]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[553] ),
        .I2(\f_permutation_l_/out_reg_n_0_[153] ),
        .I3(\out[1540]_i_4_n_0 ),
        .I4(\out[1238]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1046]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1047]_i_1 
       (.I0(\out[1558]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[554] ),
        .I2(\f_permutation_l_/out_reg_n_0_[154] ),
        .I3(\out[1541]_i_4_n_0 ),
        .I4(\out[1239]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1047]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1048]_i_1 
       (.I0(\out[1559]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[555] ),
        .I2(\f_permutation_l_/out_reg_n_0_[155] ),
        .I3(\out[1542]_i_4_n_0 ),
        .I4(\out[1240]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1048]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1049]_i_1 
       (.I0(\out[1560]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[556] ),
        .I2(\f_permutation_l_/out_reg_n_0_[156] ),
        .I3(\out[1543]_i_4_n_0 ),
        .I4(\out[1241]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1049]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[104]_i_1 
       (.I0(\out[1218]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[639] ),
        .I2(\f_permutation_l_/out_reg_n_0_[230] ),
        .I3(\out[1554]_i_3_n_0 ),
        .I4(\out[296]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1050]_i_1 
       (.I0(\out[1561]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[557] ),
        .I2(\f_permutation_l_/out_reg_n_0_[157] ),
        .I3(\out[1544]_i_4_n_0 ),
        .I4(\out[1242]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1050]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1051]_i_1 
       (.I0(\out[1562]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[558] ),
        .I2(\f_permutation_l_/out_reg_n_0_[158] ),
        .I3(\out[1545]_i_4_n_0 ),
        .I4(\out[1243]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1051]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1052]_i_1 
       (.I0(\out[1563]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[559] ),
        .I2(\f_permutation_l_/out_reg_n_0_[159] ),
        .I3(\out[1546]_i_4_n_0 ),
        .I4(\out[1244]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1052]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1053]_i_1 
       (.I0(\out[1564]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[560] ),
        .I2(\f_permutation_l_/out_reg_n_0_[160] ),
        .I3(\out[1547]_i_4_n_0 ),
        .I4(\out[1245]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1053]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1054]_i_1 
       (.I0(\out[1565]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[561] ),
        .I2(\f_permutation_l_/out_reg_n_0_[161] ),
        .I3(\out[1548]_i_4_n_0 ),
        .I4(\out[1246]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1054]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1055]_i_1 
       (.I0(\out[1566]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[562] ),
        .I2(\f_permutation_l_/out_reg_n_0_[162] ),
        .I3(\out[1549]_i_4_n_0 ),
        .I4(\out[1247]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1055]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1056]_i_1 
       (.I0(\out[1311]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[563] ),
        .I2(\f_permutation_l_/out_reg_n_0_[163] ),
        .I3(\out[1550]_i_4_n_0 ),
        .I4(\out[1248]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1056]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1057]_i_1 
       (.I0(\out[1568]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[564] ),
        .I2(\f_permutation_l_/out_reg_n_0_[164] ),
        .I3(\out[1551]_i_3_n_0 ),
        .I4(\out[1249]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1057]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1058]_i_1 
       (.I0(\out[1569]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[565] ),
        .I2(\f_permutation_l_/out_reg_n_0_[165] ),
        .I3(\out[1552]_i_4_n_0 ),
        .I4(\out[1250]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1058]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1059]_i_1 
       (.I0(\out[1570]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[566] ),
        .I2(\f_permutation_l_/out_reg_n_0_[166] ),
        .I3(\out[1553]_i_4_n_0 ),
        .I4(\out[1251]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1059]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[105]_i_1 
       (.I0(\out[1219]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[576] ),
        .I2(\f_permutation_l_/out_reg_n_0_[231] ),
        .I3(\out[1555]_i_3_n_0 ),
        .I4(\out[297]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1060]_i_1 
       (.I0(\out[1571]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[567] ),
        .I2(\f_permutation_l_/out_reg_n_0_[167] ),
        .I3(\out[1554]_i_4_n_0 ),
        .I4(\out[1252]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1060]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1061]_i_1 
       (.I0(\out[1572]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[568] ),
        .I2(\f_permutation_l_/out_reg_n_0_[168] ),
        .I3(\out[1555]_i_4_n_0 ),
        .I4(\out[1253]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1061]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1062]_i_1 
       (.I0(\out[1573]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[569] ),
        .I2(\f_permutation_l_/out_reg_n_0_[169] ),
        .I3(\out[1556]_i_4_n_0 ),
        .I4(\out[1254]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1062]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1063]_i_1 
       (.I0(\out[1574]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[570] ),
        .I2(\f_permutation_l_/out_reg_n_0_[170] ),
        .I3(\out[1557]_i_4_n_0 ),
        .I4(\out[1255]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1063]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1064]_i_1 
       (.I0(\out[1575]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[571] ),
        .I2(\f_permutation_l_/out_reg_n_0_[171] ),
        .I3(\out[1558]_i_4_n_0 ),
        .I4(\out[1256]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1064]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1065]_i_1 
       (.I0(\out[1576]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[572] ),
        .I2(\f_permutation_l_/out_reg_n_0_[172] ),
        .I3(\out[1559]_i_4_n_0 ),
        .I4(\out[1257]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1065]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1066]_i_1 
       (.I0(\out[1577]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[573] ),
        .I2(\f_permutation_l_/out_reg_n_0_[173] ),
        .I3(\out[1560]_i_4_n_0 ),
        .I4(\out[1258]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1066]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1067]_i_1 
       (.I0(\out[1578]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[574] ),
        .I2(\f_permutation_l_/out_reg_n_0_[174] ),
        .I3(\out[1561]_i_4_n_0 ),
        .I4(\out[1259]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1067]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1068]_i_1 
       (.I0(\out[1579]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[575] ),
        .I2(\f_permutation_l_/out_reg_n_0_[175] ),
        .I3(\out[1562]_i_4_n_0 ),
        .I4(\out[1260]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1068]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1069]_i_1 
       (.I0(\out[1580]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[512] ),
        .I2(\f_permutation_l_/out_reg_n_0_[176] ),
        .I3(\out[1563]_i_4_n_0 ),
        .I4(\out[1261]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1069]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[106]_i_1 
       (.I0(\out[1220]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[577] ),
        .I2(\f_permutation_l_/out_reg_n_0_[232] ),
        .I3(\out[1556]_i_3_n_0 ),
        .I4(\out[298]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[1070]_i_1 
       (.I0(\out[1581]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[513] ),
        .I2(\f_permutation_l_/out_reg_n_0_[177] ),
        .I3(\out[1564]_i_4_n_0 ),
        .I4(\out[1262]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1070]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1071]_i_1 
       (.I0(\out[1582]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[514] ),
        .I2(\f_permutation_l_/out_reg_n_0_[178] ),
        .I3(\out[1565]_i_4_n_0 ),
        .I4(\out[1263]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1071]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1072]_i_1 
       (.I0(\out[1583]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[515] ),
        .I2(\f_permutation_l_/out_reg_n_0_[179] ),
        .I3(\out[1566]_i_4_n_0 ),
        .I4(\out[1264]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1072]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1073]_i_1 
       (.I0(\out[1584]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[516] ),
        .I2(\f_permutation_l_/out_reg_n_0_[180] ),
        .I3(\out[1567]_i_3_n_0 ),
        .I4(\out[1265]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1073]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1074]_i_1 
       (.I0(\out[1585]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[517] ),
        .I2(\f_permutation_l_/out_reg_n_0_[181] ),
        .I3(\out[1568]_i_4_n_0 ),
        .I4(\out[1266]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1074]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1075]_i_1 
       (.I0(\out[1586]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[518] ),
        .I2(\f_permutation_l_/out_reg_n_0_[182] ),
        .I3(\out[1569]_i_4_n_0 ),
        .I4(\out[1267]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1075]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1076]_i_1 
       (.I0(\out[1587]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[519] ),
        .I2(\f_permutation_l_/out_reg_n_0_[183] ),
        .I3(\out[1570]_i_4_n_0 ),
        .I4(\out[1268]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1076]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1077]_i_1 
       (.I0(\out[1588]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[520] ),
        .I2(\f_permutation_l_/out_reg_n_0_[184] ),
        .I3(\out[1571]_i_4_n_0 ),
        .I4(\out[1269]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1077]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1078]_i_1 
       (.I0(\out[1589]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[521] ),
        .I2(\f_permutation_l_/out_reg_n_0_[185] ),
        .I3(\out[1572]_i_4_n_0 ),
        .I4(\out[1270]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1078]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1079]_i_1 
       (.I0(\out[1590]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[522] ),
        .I2(\f_permutation_l_/out_reg_n_0_[186] ),
        .I3(\out[1573]_i_4_n_0 ),
        .I4(\out[1271]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1079]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[107]_i_1 
       (.I0(\out[1221]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[578] ),
        .I2(\f_permutation_l_/out_reg_n_0_[233] ),
        .I3(\out[1557]_i_3_n_0 ),
        .I4(\out[299]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1080]_i_1 
       (.I0(\out[1591]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[523] ),
        .I2(\f_permutation_l_/out_reg_n_0_[187] ),
        .I3(\out[1574]_i_4_n_0 ),
        .I4(\out[1272]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1080]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1081]_i_1 
       (.I0(\out[1592]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[524] ),
        .I2(\f_permutation_l_/out_reg_n_0_[188] ),
        .I3(\out[1575]_i_4_n_0 ),
        .I4(\out[1273]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1081]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1082]_i_1 
       (.I0(\out[1593]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[525] ),
        .I2(\f_permutation_l_/out_reg_n_0_[189] ),
        .I3(\out[1576]_i_4_n_0 ),
        .I4(\out[1274]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1082]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1083]_i_1 
       (.I0(\out[1594]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[526] ),
        .I2(\f_permutation_l_/out_reg_n_0_[190] ),
        .I3(\out[1577]_i_4_n_0 ),
        .I4(\out[1275]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1083]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1084]_i_1 
       (.I0(\out[1595]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[527] ),
        .I2(\f_permutation_l_/out_reg_n_0_[191] ),
        .I3(\out[1578]_i_4_n_0 ),
        .I4(\out[1276]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1084]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1085]_i_1 
       (.I0(\out[1596]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[528] ),
        .I2(\f_permutation_l_/out_reg_n_0_[128] ),
        .I3(\out[1579]_i_4_n_0 ),
        .I4(\out[1277]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1085]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1086]_i_1 
       (.I0(\out[1597]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[529] ),
        .I2(\f_permutation_l_/out_reg_n_0_[129] ),
        .I3(\out[1580]_i_4_n_0 ),
        .I4(\out[1278]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1086]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1087]_i_1 
       (.I0(\out[1598]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[530] ),
        .I2(\f_permutation_l_/out_reg_n_0_[130] ),
        .I3(\out[1581]_i_4_n_0 ),
        .I4(\out[1279]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1087]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1088]_i_1 
       (.I0(\out[1216]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[957] ),
        .I2(\out[1088]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[131] ),
        .I4(\out[1582]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1088]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1088]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[531] ),
        .I1(\f_permutation_l_/round_in [1426]),
        .I2(\out[1599]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1555]),
        .I4(\out[1599]_i_8_n_0 ),
        .O(\out[1088]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1089]_i_1 
       (.I0(\out[1217]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[958] ),
        .I2(\out[1089]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[132] ),
        .I4(\out[1583]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1089]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1089]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[532] ),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1556]),
        .I4(\out[1536]_i_10_n_0 ),
        .O(\out[1089]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[108]_i_1 
       (.I0(\out[1539]_i_6_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[579] ),
        .I2(\f_permutation_l_/out_reg_n_0_[234] ),
        .I3(\out[1558]_i_3_n_0 ),
        .I4(\out[300]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1090]_i_1 
       (.I0(\out[1218]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[959] ),
        .I2(\out[1090]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[133] ),
        .I4(\out[1584]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1090]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1090]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[533] ),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1557]),
        .I4(\out[1537]_i_9_n_0 ),
        .O(\out[1090]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1091]_i_1 
       (.I0(\out[1219]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[896] ),
        .I2(\out[1091]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[134] ),
        .I4(\out[1585]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1091]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1091]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[534] ),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1558]),
        .I4(\out[1538]_i_6_n_0 ),
        .O(\out[1091]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1092]_i_1 
       (.I0(\out[1220]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[897] ),
        .I2(\out[1092]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[135] ),
        .I4(\out[1586]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1092]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1092]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[535] ),
        .I1(\f_permutation_l_/round_in [1430]),
        .I2(\out[1539]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1559]),
        .I4(\out[1539]_i_8_n_0 ),
        .O(\out[1092]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1093]_i_1 
       (.I0(\out[1221]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[898] ),
        .I2(\out[1093]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[136] ),
        .I4(\out[1587]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1093]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1093]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[536] ),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1560]),
        .I4(\out[1540]_i_6_n_0 ),
        .O(\out[1093]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1094]_i_1 
       (.I0(\out[1539]_i_6_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[899] ),
        .I2(\out[1094]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[137] ),
        .I4(\out[1588]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1094]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1094]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[537] ),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1561]),
        .I4(\out[1541]_i_6_n_0 ),
        .O(\out[1094]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1095]_i_1 
       (.I0(\out[1223]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[900] ),
        .I2(\out[1095]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[138] ),
        .I4(\out[1589]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1095]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1095]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[538] ),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1562]),
        .I4(\out[1542]_i_7_n_0 ),
        .O(\out[1095]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1096]_i_1 
       (.I0(\out[1224]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[901] ),
        .I2(\out[1096]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[139] ),
        .I4(\out[1590]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1096]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1096]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[539] ),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1563]),
        .I4(\out[1543]_i_10_n_0 ),
        .O(\out[1096]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1097]_i_1 
       (.I0(\out[1225]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[902] ),
        .I2(\out[1097]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[140] ),
        .I4(\out[1591]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1097]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1097]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[540] ),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1564]),
        .I4(\out[1544]_i_6_n_0 ),
        .O(\out[1097]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1098]_i_1 
       (.I0(\out[1226]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[903] ),
        .I2(\out[1098]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[141] ),
        .I4(\out[1592]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1098]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1098]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[541] ),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1565]),
        .I4(\out[1545]_i_6_n_0 ),
        .O(\out[1098]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1099]_i_1 
       (.I0(\out[1227]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[904] ),
        .I2(\out[1099]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[142] ),
        .I4(\out[1593]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1099]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1099]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[542] ),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1566]),
        .I4(\out[1546]_i_6_n_0 ),
        .O(\out[1099]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[109]_i_1 
       (.I0(\out[1223]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[580] ),
        .I2(\f_permutation_l_/out_reg_n_0_[235] ),
        .I3(\out[1559]_i_3_n_0 ),
        .I4(\out[301]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[10]_i_1 
       (.I0(\out[1588]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[200] ),
        .I2(\out[266]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1043]),
        .I4(\out[1512]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1100]_i_1 
       (.I0(\out[1228]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[905] ),
        .I2(\out[1100]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[143] ),
        .I4(\out[1594]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1100]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[543] ),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1567]),
        .I4(\out[1547]_i_6_n_0 ),
        .O(\out[1100]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1101]_i_1 
       (.I0(\out[1229]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[906] ),
        .I2(\out[1101]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[144] ),
        .I4(\out[1595]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1101]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[544] ),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1568]),
        .I4(\out[1548]_i_6_n_0 ),
        .O(\out[1101]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1102]_i_1 
       (.I0(\out[1230]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[907] ),
        .I2(\out[1102]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[145] ),
        .I4(\out[1596]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1102]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[545] ),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1569]),
        .I4(\out[1549]_i_6_n_0 ),
        .O(\out[1102]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1103]_i_1 
       (.I0(\out[1231]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[908] ),
        .I2(\out[1103]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[146] ),
        .I4(\out[1597]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1103]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[546] ),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1570]),
        .I4(\out[1550]_i_6_n_0 ),
        .O(\out[1103]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1104]_i_1 
       (.I0(\out[1232]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[909] ),
        .I2(\out[1104]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[147] ),
        .I4(\out[1598]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1104]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[547] ),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1571]),
        .I4(\out[1551]_i_9_n_0 ),
        .O(\out[1104]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1105]_i_1 
       (.I0(\out[1233]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[910] ),
        .I2(\out[1105]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[148] ),
        .I4(\out[1599]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1105]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[548] ),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1572]),
        .I4(\out[1552]_i_6_n_0 ),
        .O(\out[1105]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1106]_i_1 
       (.I0(\out[1234]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[911] ),
        .I2(\out[1106]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[149] ),
        .I4(\out[1472]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1106]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[549] ),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1573]),
        .I4(\out[1553]_i_6_n_0 ),
        .O(\out[1106]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1107]_i_1 
       (.I0(\out[1235]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[912] ),
        .I2(\out[1107]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[150] ),
        .I4(\out[1537]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1107]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[550] ),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1574]),
        .I4(\out[1554]_i_6_n_0 ),
        .O(\out[1107]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1108]_i_1 
       (.I0(\out[1236]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[913] ),
        .I2(\out[1108]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[151] ),
        .I4(\out[1538]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1108]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[551] ),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1575]),
        .I4(\out[1555]_i_6_n_0 ),
        .O(\out[1108]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1109]_i_1 
       (.I0(\out[1237]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[914] ),
        .I2(\f_permutation_l_/out_reg_n_0_[552] ),
        .I3(\out[1556]_i_3_n_0 ),
        .I4(\out[1109]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1109]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[152] ),
        .I1(\out[1539]_i_12_n_0 ),
        .I2(\f_permutation_l_/round_in [1367]),
        .I3(\f_permutation_l_/round_in [1496]),
        .I4(\out[1539]_i_14_n_0 ),
        .O(\out[1109]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[110]_i_1 
       (.I0(\out[1224]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[581] ),
        .I2(\f_permutation_l_/out_reg_n_0_[236] ),
        .I3(\out[1560]_i_3_n_0 ),
        .I4(\out[302]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1110]_i_1 
       (.I0(\out[1238]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[915] ),
        .I2(\out[1110]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[153] ),
        .I4(\out[1540]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1110]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[553] ),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1577]),
        .I4(\out[1557]_i_6_n_0 ),
        .O(\out[1110]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1111]_i_1 
       (.I0(\out[1239]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[916] ),
        .I2(\out[1111]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[154] ),
        .I4(\out[1541]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1111]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[554] ),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1578]),
        .I4(\out[1558]_i_6_n_0 ),
        .O(\out[1111]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1112]_i_1 
       (.I0(\out[1240]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[917] ),
        .I2(\out[1112]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[155] ),
        .I4(\out[1542]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1112]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[555] ),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1579]),
        .I4(\out[1559]_i_6_n_0 ),
        .O(\out[1112]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1113]_i_1 
       (.I0(\out[1241]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[918] ),
        .I2(\out[1113]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[156] ),
        .I4(\out[1543]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1113]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[556] ),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1580]),
        .I4(\out[1560]_i_6_n_0 ),
        .O(\out[1113]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1114]_i_1 
       (.I0(\out[1242]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[919] ),
        .I2(\out[1114]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[157] ),
        .I4(\out[1544]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1114]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[557] ),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1581]),
        .I4(\out[1561]_i_6_n_0 ),
        .O(\out[1114]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1115]_i_1 
       (.I0(\out[1243]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[920] ),
        .I2(\out[1115]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[158] ),
        .I4(\out[1545]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1115]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[558] ),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1582]),
        .I4(\out[1562]_i_6_n_0 ),
        .O(\out[1115]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1116]_i_1 
       (.I0(\out[1244]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[921] ),
        .I2(\out[1116]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[159] ),
        .I4(\out[1546]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1116]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[559] ),
        .I1(\f_permutation_l_/round_in [1454]),
        .I2(\out[1563]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1583]),
        .I4(\out[1563]_i_6_n_0 ),
        .O(\out[1116]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1117]_i_1 
       (.I0(\out[1245]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[922] ),
        .I2(\out[1117]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[160] ),
        .I4(\out[1547]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1117]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[560] ),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1584]),
        .I4(\out[1564]_i_6_n_0 ),
        .O(\out[1117]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1118]_i_1 
       (.I0(\out[1246]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[923] ),
        .I2(\out[1118]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[161] ),
        .I4(\out[1548]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1118]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[561] ),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1585]),
        .I4(\out[1565]_i_6_n_0 ),
        .O(\out[1118]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1119]_i_1 
       (.I0(\out[1247]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[924] ),
        .I2(\out[1119]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[162] ),
        .I4(\out[1549]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1119]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[562] ),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1586]),
        .I4(\out[1566]_i_6_n_0 ),
        .O(\out[1119]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[111]_i_1 
       (.I0(\out[1225]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[582] ),
        .I2(\f_permutation_l_/out_reg_n_0_[237] ),
        .I3(\out[1561]_i_3_n_0 ),
        .I4(\out[303]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1120]_i_1 
       (.I0(\out[1248]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[925] ),
        .I2(\out[1120]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[163] ),
        .I4(\out[1550]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1120]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[563] ),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1587]),
        .I4(\out[1567]_i_9_n_0 ),
        .O(\out[1120]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1121]_i_1 
       (.I0(\out[1249]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[926] ),
        .I2(\out[1121]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[164] ),
        .I4(\out[1551]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1121]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[564] ),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1588]),
        .I4(\out[1568]_i_6_n_0 ),
        .O(\out[1121]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1122]_i_1 
       (.I0(\out[1250]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[927] ),
        .I2(\out[1122]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[165] ),
        .I4(\out[1552]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1122]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[565] ),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1589]),
        .I4(\out[1569]_i_6_n_0 ),
        .O(\out[1122]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1123]_i_1 
       (.I0(\out[1251]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[928] ),
        .I2(\out[1123]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[166] ),
        .I4(\out[1553]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1123]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[566] ),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1590]),
        .I4(\out[1570]_i_6_n_0 ),
        .O(\out[1123]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1124]_i_1 
       (.I0(\out[1252]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[929] ),
        .I2(\out[1124]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[167] ),
        .I4(\out[1554]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1124]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[567] ),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1591]),
        .I4(\out[1571]_i_6_n_0 ),
        .O(\out[1124]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1125]_i_1 
       (.I0(\out[1253]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[930] ),
        .I2(\out[1125]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[168] ),
        .I4(\out[1555]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1125]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[568] ),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1592]),
        .I4(\out[1572]_i_6_n_0 ),
        .O(\out[1125]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1126]_i_1 
       (.I0(\out[1254]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[931] ),
        .I2(\out[1126]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[169] ),
        .I4(\out[1556]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1126]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[569] ),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1593]),
        .I4(\out[1573]_i_6_n_0 ),
        .O(\out[1126]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1127]_i_1 
       (.I0(\out[1255]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[932] ),
        .I2(\out[1127]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[170] ),
        .I4(\out[1557]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1127]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[570] ),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1594]),
        .I4(\out[1574]_i_6_n_0 ),
        .O(\out[1127]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1128]_i_1 
       (.I0(\out[1256]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[933] ),
        .I2(\out[1128]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[171] ),
        .I4(\out[1558]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1128]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1128]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[571] ),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1595]),
        .I4(\out[1575]_i_6_n_0 ),
        .O(\out[1128]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1129]_i_1 
       (.I0(\out[1257]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[934] ),
        .I2(\out[1129]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[172] ),
        .I4(\out[1559]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1129]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1129]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[572] ),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1596]),
        .I4(\out[1576]_i_6_n_0 ),
        .O(\out[1129]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[112]_i_1 
       (.I0(\out[1226]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[583] ),
        .I2(\f_permutation_l_/out_reg_n_0_[238] ),
        .I3(\out[1562]_i_3_n_0 ),
        .I4(\out[304]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1130]_i_1 
       (.I0(\out[1258]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[935] ),
        .I2(\out[1130]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[173] ),
        .I4(\out[1560]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1130]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1130]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[573] ),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1597]),
        .I4(\out[1577]_i_6_n_0 ),
        .O(\out[1130]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1131]_i_1 
       (.I0(\out[1259]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[936] ),
        .I2(\out[1131]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[174] ),
        .I4(\out[1561]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1131]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1131]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[574] ),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1598]),
        .I4(\out[1578]_i_6_n_0 ),
        .O(\out[1131]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1132]_i_1 
       (.I0(\out[1260]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[937] ),
        .I2(\out[1132]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[175] ),
        .I4(\out[1562]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1132]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1132]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[575] ),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1599]),
        .I4(\out[1579]_i_7_n_0 ),
        .O(\out[1132]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1133]_i_1 
       (.I0(\out[1261]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[938] ),
        .I2(\out[1133]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[176] ),
        .I4(\out[1563]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1133]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1133]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[512] ),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1536]),
        .I4(\out[1580]_i_6_n_0 ),
        .O(\out[1133]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1134]_i_1 
       (.I0(\out[1262]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[939] ),
        .I2(\out[1134]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[177] ),
        .I4(\out[1564]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1134]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1134]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[513] ),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1537]),
        .I4(\out[1581]_i_6_n_0 ),
        .O(\out[1134]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1135]_i_1 
       (.I0(\out[1263]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[940] ),
        .I2(\out[1135]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[178] ),
        .I4(\out[1565]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1135]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1135]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[514] ),
        .I1(\f_permutation_l_/round_in [1409]),
        .I2(\out[1582]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1538]),
        .I4(\out[1582]_i_6_n_0 ),
        .O(\out[1135]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1136]_i_1 
       (.I0(\out[1264]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[941] ),
        .I2(\out[1136]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[179] ),
        .I4(\out[1566]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1136]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1136]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[515] ),
        .I1(\f_permutation_l_/round_in [1410]),
        .I2(\out[1583]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1539]),
        .I4(\out[1583]_i_6_n_0 ),
        .O(\out[1136]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1137]_i_1 
       (.I0(\out[1265]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[942] ),
        .I2(\out[1137]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[180] ),
        .I4(\out[1567]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1137]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1137]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[516] ),
        .I1(\f_permutation_l_/round_in [1411]),
        .I2(\out[1584]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1540]),
        .I4(\out[1584]_i_6_n_0 ),
        .O(\out[1137]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1138]_i_1 
       (.I0(\out[1266]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[943] ),
        .I2(\out[1138]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[181] ),
        .I4(\out[1568]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1138]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1138]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[517] ),
        .I1(\f_permutation_l_/round_in [1412]),
        .I2(\out[1585]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1541]),
        .I4(\out[1585]_i_6_n_0 ),
        .O(\out[1138]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1139]_i_1 
       (.I0(\out[1267]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[944] ),
        .I2(\out[1139]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[182] ),
        .I4(\out[1569]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1139]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1139]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[518] ),
        .I1(\f_permutation_l_/round_in [1413]),
        .I2(\out[1586]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1542]),
        .I4(\out[1586]_i_6_n_0 ),
        .O(\out[1139]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[113]_i_1 
       (.I0(\out[1227]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[584] ),
        .I2(\f_permutation_l_/out_reg_n_0_[239] ),
        .I3(\out[1563]_i_3_n_0 ),
        .I4(\out[305]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1140]_i_1 
       (.I0(\out[1268]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[945] ),
        .I2(\out[1140]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[183] ),
        .I4(\out[1570]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1140]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1140]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[519] ),
        .I1(\f_permutation_l_/round_in [1414]),
        .I2(\out[1587]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1543]),
        .I4(\out[1587]_i_6_n_0 ),
        .O(\out[1140]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1141]_i_1 
       (.I0(\out[1269]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[946] ),
        .I2(\out[1141]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[184] ),
        .I4(\out[1571]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1141]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1141]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[520] ),
        .I1(\f_permutation_l_/round_in [1415]),
        .I2(\out[1588]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1544]),
        .I4(\out[1588]_i_6_n_0 ),
        .O(\out[1141]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1142]_i_1 
       (.I0(\out[1270]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[947] ),
        .I2(\out[1142]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[185] ),
        .I4(\out[1572]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1142]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1142]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[521] ),
        .I1(\f_permutation_l_/round_in [1416]),
        .I2(\out[1589]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1545]),
        .I4(\out[1589]_i_6_n_0 ),
        .O(\out[1142]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1143]_i_1 
       (.I0(\out[1271]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[948] ),
        .I2(\out[1143]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[186] ),
        .I4(\out[1573]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1143]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1143]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[522] ),
        .I1(\f_permutation_l_/round_in [1417]),
        .I2(\out[1590]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1546]),
        .I4(\out[1590]_i_6_n_0 ),
        .O(\out[1143]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1144]_i_1 
       (.I0(\out[1272]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[949] ),
        .I2(\out[1144]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[187] ),
        .I4(\out[1574]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1144]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1144]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[523] ),
        .I1(\f_permutation_l_/round_in [1418]),
        .I2(\out[1591]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1547]),
        .I4(\out[1591]_i_6_n_0 ),
        .O(\out[1144]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1145]_i_1 
       (.I0(\out[1273]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[950] ),
        .I2(\out[1145]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[188] ),
        .I4(\out[1575]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1145]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1145]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[524] ),
        .I1(\f_permutation_l_/round_in [1419]),
        .I2(\out[1592]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1548]),
        .I4(\out[1592]_i_6_n_0 ),
        .O(\out[1145]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1146]_i_1 
       (.I0(\out[1274]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[951] ),
        .I2(\out[1146]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[189] ),
        .I4(\out[1576]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1146]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1146]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[525] ),
        .I1(\f_permutation_l_/round_in [1420]),
        .I2(\out[1593]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1549]),
        .I4(\out[1593]_i_6_n_0 ),
        .O(\out[1146]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1147]_i_1 
       (.I0(\out[1275]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[952] ),
        .I2(\out[1147]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[190] ),
        .I4(\out[1577]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1147]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1147]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[526] ),
        .I1(\f_permutation_l_/round_in [1421]),
        .I2(\out[1594]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1550]),
        .I4(\out[1594]_i_6_n_0 ),
        .O(\out[1147]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1148]_i_1 
       (.I0(\out[1276]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[953] ),
        .I2(\out[1148]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[191] ),
        .I4(\out[1578]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1148]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1148]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[527] ),
        .I1(\f_permutation_l_/round_in [1422]),
        .I2(\out[1595]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1551]),
        .I4(\out[1595]_i_6_n_0 ),
        .O(\out[1148]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1149]_i_1 
       (.I0(\out[1277]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[954] ),
        .I2(\out[1149]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[128] ),
        .I4(\out[1579]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1149]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1149]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[528] ),
        .I1(\f_permutation_l_/round_in [1423]),
        .I2(\out[1596]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1552]),
        .I4(\out[1596]_i_6_n_0 ),
        .O(\out[1149]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[114]_i_1 
       (.I0(\out[1228]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[585] ),
        .I2(\f_permutation_l_/out_reg_n_0_[240] ),
        .I3(\out[1564]_i_3_n_0 ),
        .I4(\out[306]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1150]_i_1 
       (.I0(\out[1278]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[955] ),
        .I2(\out[1150]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[129] ),
        .I4(\out[1580]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1150]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1150]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[529] ),
        .I1(\f_permutation_l_/round_in [1424]),
        .I2(\out[1597]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1553]),
        .I4(\out[1597]_i_6_n_0 ),
        .O(\out[1150]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1151]_i_1 
       (.I0(\out[1279]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[956] ),
        .I2(\out[1151]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[130] ),
        .I4(\out[1581]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1151]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1151]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[530] ),
        .I1(\f_permutation_l_/round_in [1425]),
        .I2(\out[1598]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1554]),
        .I4(\out[1598]_i_6_n_0 ),
        .O(\out[1151]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1152]_i_1 
       (.I0(\out[1466]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1004] ),
        .I2(\out[1152]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[531] ),
        .I4(\out[1343]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1152]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1152]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[957] ),
        .I1(\f_permutation_l_/round_in [1532]),
        .I2(\out[1575]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[1152]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1153]_i_1 
       (.I0(\out[1467]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1005] ),
        .I2(\out[1153]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[532] ),
        .I4(\out[1280]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1153]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1153]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[958] ),
        .I1(\f_permutation_l_/round_in [1533]),
        .I2(\out[1576]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[1153]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1154]_i_1 
       (.I0(\out[1468]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1006] ),
        .I2(\out[1154]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[533] ),
        .I4(\out[1281]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1154]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1154]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[959] ),
        .I1(\f_permutation_l_/round_in [1534]),
        .I2(\out[1577]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[1154]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1155]_i_1 
       (.I0(\out[1469]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1007] ),
        .I2(\out[1155]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[534] ),
        .I4(\out[1538]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1155]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1155]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[896] ),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[1155]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1156]_i_1 
       (.I0(\out[1470]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1008] ),
        .I2(\out[1156]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[535] ),
        .I4(\out[1539]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1156]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1156]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[897] ),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[1156]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1157]_i_1 
       (.I0(\out[1471]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1009] ),
        .I2(\out[1157]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[536] ),
        .I4(\out[1540]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1157]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1157]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[898] ),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[1157]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1158]_i_1 
       (.I0(\out[1408]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1010] ),
        .I2(\out[1158]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[537] ),
        .I4(\out[1541]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1158]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1158]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[899] ),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[1158]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1159]_i_1 
       (.I0(\out[1409]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1011] ),
        .I2(\out[1159]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[538] ),
        .I4(\out[1542]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1159]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1159]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[900] ),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[1159]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[115]_i_1 
       (.I0(\out[1229]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[586] ),
        .I2(\f_permutation_l_/out_reg_n_0_[241] ),
        .I3(\out[1565]_i_3_n_0 ),
        .I4(\out[307]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1160]_i_1 
       (.I0(\out[1410]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1012] ),
        .I2(\out[1160]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[539] ),
        .I4(\out[1287]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1160]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1160]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[901] ),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[1160]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1161]_i_1 
       (.I0(\out[1411]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1013] ),
        .I2(\out[1161]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[540] ),
        .I4(\out[1544]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1161]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1161]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[902] ),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[1161]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1162]_i_1 
       (.I0(\out[1412]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1014] ),
        .I2(\out[1162]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[541] ),
        .I4(\out[1545]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1162]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1162]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[903] ),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[1162]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1163]_i_1 
       (.I0(\out[1413]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1015] ),
        .I2(\out[1163]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[542] ),
        .I4(\out[1546]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1163]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1163]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[904] ),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[1163]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1164]_i_1 
       (.I0(\out[1414]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1016] ),
        .I2(\out[1164]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[543] ),
        .I4(\out[1547]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1164]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1164]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[905] ),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[1164]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1165]_i_1 
       (.I0(\out[1415]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1017] ),
        .I2(\out[1165]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[544] ),
        .I4(\out[1548]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1165]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1165]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[906] ),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[1165]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1166]_i_1 
       (.I0(\out[1416]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1018] ),
        .I2(\out[1166]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[545] ),
        .I4(\out[1549]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1166]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1166]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[907] ),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[1166]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1167]_i_1 
       (.I0(\out[1417]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1019] ),
        .I2(\out[1167]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[546] ),
        .I4(\out[1550]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1167]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1167]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[908] ),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[1167]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1168]_i_1 
       (.I0(\out[1418]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1020] ),
        .I2(\out[1168]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[547] ),
        .I4(\out[1295]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1168]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1168]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[909] ),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[1168]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1169]_i_1 
       (.I0(\out[1419]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1021] ),
        .I2(\out[1169]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[548] ),
        .I4(\out[1552]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1169]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1169]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[910] ),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[1169]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[116]_i_1 
       (.I0(\out[1230]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[587] ),
        .I2(\f_permutation_l_/out_reg_n_0_[242] ),
        .I3(\out[1566]_i_3_n_0 ),
        .I4(\out[308]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1170]_i_1 
       (.I0(\out[1420]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1022] ),
        .I2(\out[1170]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[549] ),
        .I4(\out[1553]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1170]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1170]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[911] ),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[1170]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1171]_i_1 
       (.I0(\out[1421]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1023] ),
        .I2(\out[1171]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[550] ),
        .I4(\out[1554]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1171]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1171]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[912] ),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[1171]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1172]_i_1 
       (.I0(\out[1422]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[960] ),
        .I2(\out[1172]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[551] ),
        .I4(\out[1555]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1172]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1172]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[913] ),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[1172]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1173]_i_1 
       (.I0(\out[1423]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[961] ),
        .I2(\out[1173]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[552] ),
        .I4(\out[1556]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1173]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1173]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[914] ),
        .I1(\f_permutation_l_/round_in [1298]),
        .I2(\out[1554]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[1173]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1174]_i_1 
       (.I0(\out[1424]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[962] ),
        .I2(\out[1174]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[553] ),
        .I4(\out[1557]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1174]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1174]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[915] ),
        .I1(\f_permutation_l_/round_in [1299]),
        .I2(\out[1555]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[1174]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1175]_i_1 
       (.I0(\out[1425]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[963] ),
        .I2(\out[1175]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[554] ),
        .I4(\out[1558]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1175]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1175]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[916] ),
        .I1(\f_permutation_l_/round_in [1300]),
        .I2(\out[1556]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[1175]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1176]_i_1 
       (.I0(\out[1426]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[964] ),
        .I2(\out[1176]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[555] ),
        .I4(\out[1559]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1176]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1176]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[917] ),
        .I1(\f_permutation_l_/round_in [1301]),
        .I2(\out[1557]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[1176]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1177]_i_1 
       (.I0(\out[1427]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[965] ),
        .I2(\out[1177]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[556] ),
        .I4(\out[1560]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1177]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1177]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[918] ),
        .I1(\out[1536]_i_14_n_0 ),
        .I2(\f_permutation_l_/round_in [1493]),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[1177]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1178]_i_1 
       (.I0(\out[1428]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[966] ),
        .I2(\out[1178]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[557] ),
        .I4(\out[1561]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1178]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1178]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[919] ),
        .I1(\f_permutation_l_/round_in [1494]),
        .I2(\out[1537]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[1178]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1179]_i_1 
       (.I0(\out[1429]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[967] ),
        .I2(\out[1179]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[558] ),
        .I4(\out[1562]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1179]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1179]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[920] ),
        .I1(\f_permutation_l_/round_in [1495]),
        .I2(\out[1538]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[1179]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[117]_i_1 
       (.I0(\out[1231]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[588] ),
        .I2(\f_permutation_l_/out_reg_n_0_[243] ),
        .I3(\out[1311]_i_3_n_0 ),
        .I4(\out[309]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1180]_i_1 
       (.I0(\out[1430]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[968] ),
        .I2(\out[1180]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[559] ),
        .I4(\out[1563]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1180]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1180]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[921] ),
        .I1(\f_permutation_l_/round_in [1496]),
        .I2(\out[1539]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[1180]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1181]_i_1 
       (.I0(\out[1431]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[969] ),
        .I2(\out[1181]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[560] ),
        .I4(\out[1564]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1181]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1181]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[922] ),
        .I1(\f_permutation_l_/round_in [1497]),
        .I2(\out[1540]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[1181]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1182]_i_1 
       (.I0(\out[1432]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[970] ),
        .I2(\out[1182]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[561] ),
        .I4(\out[1565]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1182]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1182]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[923] ),
        .I1(\f_permutation_l_/round_in [1498]),
        .I2(\out[1541]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[1182]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1183]_i_1 
       (.I0(\out[1433]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[971] ),
        .I2(\out[1183]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[562] ),
        .I4(\out[1566]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1183]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1183]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[924] ),
        .I1(\f_permutation_l_/round_in [1499]),
        .I2(\out[1542]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[1183]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1184]_i_1 
       (.I0(\out[1434]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[972] ),
        .I2(\out[1184]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[563] ),
        .I4(\out[1311]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1184]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1184]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[925] ),
        .I1(\f_permutation_l_/round_in [1500]),
        .I2(\out[1543]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[1184]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1185]_i_1 
       (.I0(\out[1435]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[973] ),
        .I2(\out[1185]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[564] ),
        .I4(\out[1568]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1185]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1185]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[926] ),
        .I1(\f_permutation_l_/round_in [1501]),
        .I2(\out[1544]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[1185]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1186]_i_1 
       (.I0(\out[1436]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[974] ),
        .I2(\out[1186]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[565] ),
        .I4(\out[1569]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1186]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1186]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[927] ),
        .I1(\f_permutation_l_/round_in [1502]),
        .I2(\out[1545]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[1186]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1187]_i_1 
       (.I0(\out[1437]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[975] ),
        .I2(\out[1187]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[566] ),
        .I4(\out[1570]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1187]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1187]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[928] ),
        .I1(\f_permutation_l_/round_in [1503]),
        .I2(\out[1546]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[1187]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1188]_i_1 
       (.I0(\out[1438]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[976] ),
        .I2(\out[1188]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[567] ),
        .I4(\out[1571]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1188]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1188]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[929] ),
        .I1(\f_permutation_l_/round_in [1504]),
        .I2(\out[1547]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[1188]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1189]_i_1 
       (.I0(\out[1439]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[977] ),
        .I2(\out[1189]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[568] ),
        .I4(\out[1572]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1189]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1189]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[930] ),
        .I1(\f_permutation_l_/round_in [1505]),
        .I2(\out[1548]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[1189]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[118]_i_1 
       (.I0(\out[1232]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[589] ),
        .I2(\f_permutation_l_/out_reg_n_0_[244] ),
        .I3(\out[1568]_i_3_n_0 ),
        .I4(\out[310]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1190]_i_1 
       (.I0(\out[1440]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[978] ),
        .I2(\out[1190]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[569] ),
        .I4(\out[1573]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1190]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1190]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[931] ),
        .I1(\f_permutation_l_/round_in [1506]),
        .I2(\out[1549]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[1190]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1191]_i_1 
       (.I0(\out[1441]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[979] ),
        .I2(\out[1191]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[570] ),
        .I4(\out[1574]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1191]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1191]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[932] ),
        .I1(\f_permutation_l_/round_in [1507]),
        .I2(\out[1550]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[1191]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1192]_i_1 
       (.I0(\out[1442]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[980] ),
        .I2(\out[1192]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[571] ),
        .I4(\out[1575]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1192]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1192]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[933] ),
        .I1(\f_permutation_l_/round_in [1508]),
        .I2(\out[1551]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[1192]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1193]_i_1 
       (.I0(\out[1443]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[981] ),
        .I2(\out[1193]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[572] ),
        .I4(\out[1576]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1193]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1193]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[934] ),
        .I1(\f_permutation_l_/round_in [1509]),
        .I2(\out[1552]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[1193]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1194]_i_1 
       (.I0(\out[1444]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[982] ),
        .I2(\out[1194]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[573] ),
        .I4(\out[1577]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1194]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1194]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[935] ),
        .I1(\f_permutation_l_/round_in [1510]),
        .I2(\out[1553]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[1194]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1195]_i_1 
       (.I0(\out[1445]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[983] ),
        .I2(\out[1195]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[574] ),
        .I4(\out[1578]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1195]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1195]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[936] ),
        .I1(\f_permutation_l_/round_in [1511]),
        .I2(\out[1554]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[1195]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1196]_i_1 
       (.I0(\out[1446]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[984] ),
        .I2(\out[1196]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[575] ),
        .I4(\out[1579]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1196]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1196]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[937] ),
        .I1(\f_permutation_l_/round_in [1512]),
        .I2(\out[1555]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[1196]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1197]_i_1 
       (.I0(\out[1447]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[985] ),
        .I2(\out[1197]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[512] ),
        .I4(\out[1580]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1197]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1197]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[938] ),
        .I1(\f_permutation_l_/round_in [1513]),
        .I2(\out[1556]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[1197]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1198]_i_1 
       (.I0(\out[1448]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[986] ),
        .I2(\out[1198]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[513] ),
        .I4(\out[1581]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1198]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1198]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[939] ),
        .I1(\f_permutation_l_/round_in [1514]),
        .I2(\out[1557]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[1198]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1199]_i_1 
       (.I0(\out[1449]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[987] ),
        .I2(\out[1199]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[514] ),
        .I4(\out[1582]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1199]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1199]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[940] ),
        .I1(\f_permutation_l_/round_in [1515]),
        .I2(\out[1558]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[1199]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[119]_i_1 
       (.I0(\out[1233]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[590] ),
        .I2(\f_permutation_l_/out_reg_n_0_[245] ),
        .I3(\out[1569]_i_3_n_0 ),
        .I4(\out[311]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[11]_i_1 
       (.I0(\out[1589]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[201] ),
        .I2(\out[267]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1044]),
        .I4(\out[1513]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1200]_i_1 
       (.I0(\out[1450]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[988] ),
        .I2(\out[1200]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[515] ),
        .I4(\out[1583]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1200]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1200]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[941] ),
        .I1(\f_permutation_l_/round_in [1516]),
        .I2(\out[1559]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[1200]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1201]_i_1 
       (.I0(\out[1451]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[989] ),
        .I2(\out[1201]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[516] ),
        .I4(\out[1584]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1201]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1201]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[942] ),
        .I1(\f_permutation_l_/round_in [1517]),
        .I2(\out[1560]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[1201]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1202]_i_1 
       (.I0(\out[1452]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[990] ),
        .I2(\out[1202]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[517] ),
        .I4(\out[1585]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1202]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1202]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[943] ),
        .I1(\f_permutation_l_/round_in [1518]),
        .I2(\out[1561]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[1202]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1203]_i_1 
       (.I0(\out[1453]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[991] ),
        .I2(\out[1203]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[518] ),
        .I4(\out[1586]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1203]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1203]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[944] ),
        .I1(\f_permutation_l_/round_in [1519]),
        .I2(\out[1562]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[1203]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1204]_i_1 
       (.I0(\out[1454]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[992] ),
        .I2(\out[1204]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[519] ),
        .I4(\out[1587]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1204]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1204]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[945] ),
        .I1(\f_permutation_l_/round_in [1520]),
        .I2(\out[1563]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[1204]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1205]_i_1 
       (.I0(\out[1455]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[993] ),
        .I2(\out[1205]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[520] ),
        .I4(\out[1588]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1205]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1205]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[946] ),
        .I1(\f_permutation_l_/round_in [1521]),
        .I2(\out[1564]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[1205]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1206]_i_1 
       (.I0(\out[1456]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[994] ),
        .I2(\out[1206]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[521] ),
        .I4(\out[1589]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1206]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1206]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[947] ),
        .I1(\f_permutation_l_/round_in [1522]),
        .I2(\out[1565]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[1206]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1207]_i_1 
       (.I0(\out[1457]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[995] ),
        .I2(\out[1207]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[522] ),
        .I4(\out[1590]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1207]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1207]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[948] ),
        .I1(\f_permutation_l_/round_in [1523]),
        .I2(\out[1566]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[1207]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1208]_i_1 
       (.I0(\out[1458]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[996] ),
        .I2(\out[1208]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[523] ),
        .I4(\out[1591]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1208]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1208]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[949] ),
        .I1(\f_permutation_l_/round_in [1524]),
        .I2(\out[1567]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[1208]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1209]_i_1 
       (.I0(\out[1459]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[997] ),
        .I2(\out[1209]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[524] ),
        .I4(\out[1592]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1209]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1209]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[950] ),
        .I1(\f_permutation_l_/round_in [1525]),
        .I2(\out[1568]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[1209]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[120]_i_1 
       (.I0(\out[1234]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[591] ),
        .I2(\f_permutation_l_/out_reg_n_0_[246] ),
        .I3(\out[1570]_i_3_n_0 ),
        .I4(\out[312]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1210]_i_1 
       (.I0(\out[1460]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[998] ),
        .I2(\out[1210]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[525] ),
        .I4(\out[1593]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1210]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1210]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[951] ),
        .I1(\f_permutation_l_/round_in [1526]),
        .I2(\out[1569]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[1210]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1211]_i_1 
       (.I0(\out[1461]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[999] ),
        .I2(\out[1211]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[526] ),
        .I4(\out[1594]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1211]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1211]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[952] ),
        .I1(\f_permutation_l_/round_in [1527]),
        .I2(\out[1570]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[1211]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1212]_i_1 
       (.I0(\out[1462]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1000] ),
        .I2(\out[1212]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[527] ),
        .I4(\out[1595]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1212]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1212]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[953] ),
        .I1(\f_permutation_l_/round_in [1528]),
        .I2(\out[1571]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[1212]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1213]_i_1 
       (.I0(\out[1463]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1001] ),
        .I2(\out[1213]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[528] ),
        .I4(\out[1596]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1213]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1213]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[954] ),
        .I1(\f_permutation_l_/round_in [1529]),
        .I2(\out[1572]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[1213]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1214]_i_1 
       (.I0(\out[1464]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1002] ),
        .I2(\out[1214]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[529] ),
        .I4(\out[1597]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1214]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1214]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[955] ),
        .I1(\f_permutation_l_/round_in [1530]),
        .I2(\out[1573]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[1214]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1215]_i_1 
       (.I0(\out[1465]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1003] ),
        .I2(\out[1215]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[530] ),
        .I4(\out[1598]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1215]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1215]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[956] ),
        .I1(\f_permutation_l_/round_in [1531]),
        .I2(\out[1574]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[1215]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1216]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1004] ),
        .I1(\out[1466]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[957] ),
        .I3(\out[1216]_i_2_n_0 ),
        .I4(\out[1216]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1216]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1216]_i_2 
       (.I0(\out[1597]_i_14_n_0 ),
        .I1(padder_out_1[261]),
        .I2(out[197]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1575]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1532]),
        .O(\out[1216]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1216]_i_3 
       (.I0(\f_permutation_l_/round_in [1380]),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[1216]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1217]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1005] ),
        .I1(\out[1467]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[958] ),
        .I3(\out[1217]_i_2_n_0 ),
        .I4(\out[1217]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1217]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1217]_i_2 
       (.I0(\out[1598]_i_14_n_0 ),
        .I1(padder_out_1[262]),
        .I2(out[198]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1576]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1533]),
        .O(\out[1217]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1217]_i_3 
       (.I0(\f_permutation_l_/round_in [1381]),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[1217]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1218]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1006] ),
        .I1(\out[1468]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[959] ),
        .I3(\out[1218]_i_2_n_0 ),
        .I4(\out[1218]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1218]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1218]_i_2 
       (.I0(\out[1599]_i_14_n_0 ),
        .I1(padder_out_1[263]),
        .I2(out[199]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1577]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1534]),
        .O(\out[1218]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1218]_i_3 
       (.I0(\f_permutation_l_/round_in [1382]),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[1218]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1219]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1007] ),
        .I1(\out[1469]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[896] ),
        .I3(\out[1219]_i_2_n_0 ),
        .I4(\out[1219]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1219]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1219]_i_2 
       (.I0(\out[1536]_i_19_n_0 ),
        .I1(padder_out_1[455]),
        .I2(out[391]),
        .I3(\i[0]_i_1__0_n_0 ),
        .I4(\out[1536]_i_17_n_0 ),
        .I5(\f_permutation_l_/round_in [1280]),
        .O(\out[1219]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1219]_i_3 
       (.I0(\f_permutation_l_/round_in [1383]),
        .I1(\f_permutation_l_/round_in [1447]),
        .I2(\out[1556]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[1219]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[121]_i_1 
       (.I0(\out[1235]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[592] ),
        .I2(\f_permutation_l_/out_reg_n_0_[247] ),
        .I3(\out[1571]_i_3_n_0 ),
        .I4(\out[313]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1220]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1008] ),
        .I1(\out[1470]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[897] ),
        .I3(\out[1220]_i_2_n_0 ),
        .I4(\out[1220]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1220]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1220]_i_2 
       (.I0(\out[1537]_i_17_n_0 ),
        .I1(padder_out_1[504]),
        .I2(out[440]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1537]_i_15_n_0 ),
        .I5(\f_permutation_l_/round_in [1281]),
        .O(\out[1220]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1220]_i_3 
       (.I0(\f_permutation_l_/round_in [1384]),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[1220]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1221]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1009] ),
        .I1(\out[1471]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[898] ),
        .I3(\out[1221]_i_2_n_0 ),
        .I4(\out[1221]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1221]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1221]_i_2 
       (.I0(\out[1538]_i_16_n_0 ),
        .I1(padder_out_1[505]),
        .I2(out[441]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1538]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1282]),
        .O(\out[1221]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1221]_i_3 
       (.I0(\f_permutation_l_/round_in [1385]),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[1221]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1222]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1010] ),
        .I1(\out[1408]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[899] ),
        .I3(\out[1539]_i_6_n_0 ),
        .I4(\out[1222]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1222]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1222]_i_2 
       (.I0(\f_permutation_l_/round_in [1386]),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[1222]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1223]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1011] ),
        .I1(\out[1409]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[900] ),
        .I3(\out[1223]_i_2_n_0 ),
        .I4(\out[1223]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1223]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1223]_i_2 
       (.I0(\out[1540]_i_16_n_0 ),
        .I1(padder_out_1[507]),
        .I2(out[443]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1540]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1284]),
        .O(\out[1223]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1223]_i_3 
       (.I0(\f_permutation_l_/round_in [1387]),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[1223]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1224]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1012] ),
        .I1(\out[1410]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[901] ),
        .I3(\out[1224]_i_2_n_0 ),
        .I4(\out[1224]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1224]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1224]_i_2 
       (.I0(\out[1541]_i_16_n_0 ),
        .I1(padder_out_1[508]),
        .I2(out[444]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1541]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1285]),
        .O(\out[1224]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1224]_i_3 
       (.I0(\f_permutation_l_/round_in [1388]),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[1224]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1225]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1013] ),
        .I1(\out[1411]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[902] ),
        .I3(\out[1225]_i_2_n_0 ),
        .I4(\out[1225]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1225]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1225]_i_2 
       (.I0(\out[1542]_i_18_n_0 ),
        .I1(padder_out_1[509]),
        .I2(out[445]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1542]_i_16_n_0 ),
        .I5(\f_permutation_l_/round_in [1286]),
        .O(\out[1225]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1225]_i_3 
       (.I0(\f_permutation_l_/round_in [1389]),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[1225]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1226]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1014] ),
        .I1(\out[1412]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[903] ),
        .I3(\out[1226]_i_2_n_0 ),
        .I4(\out[1226]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1226]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1226]_i_2 
       (.I0(\out[1543]_i_19_n_0 ),
        .I1(padder_out_1[510]),
        .I2(out[446]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1543]_i_17_n_0 ),
        .I5(\f_permutation_l_/round_in [1287]),
        .O(\out[1226]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1226]_i_3 
       (.I0(\f_permutation_l_/round_in [1390]),
        .I1(\f_permutation_l_/round_in [1454]),
        .I2(\out[1563]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[1226]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1227]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1015] ),
        .I1(\out[1413]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[904] ),
        .I3(\out[1227]_i_2_n_0 ),
        .I4(\out[1227]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1227]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1227]_i_2 
       (.I0(\out[1544]_i_16_n_0 ),
        .I1(padder_out_1[511]),
        .I2(out[447]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1544]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1288]),
        .O(\out[1227]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1227]_i_3 
       (.I0(\f_permutation_l_/round_in [1391]),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[1227]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1228]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1016] ),
        .I1(\out[1414]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[905] ),
        .I3(\out[1228]_i_2_n_0 ),
        .I4(\out[1228]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1228]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1228]_i_2 
       (.I0(\out[1545]_i_16_n_0 ),
        .I1(padder_out_1[496]),
        .I2(out[432]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1545]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1289]),
        .O(\out[1228]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1228]_i_3 
       (.I0(\f_permutation_l_/round_in [1392]),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[1228]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1229]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1017] ),
        .I1(\out[1415]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[906] ),
        .I3(\out[1229]_i_2_n_0 ),
        .I4(\out[1229]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1229]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1229]_i_2 
       (.I0(\out[1546]_i_16_n_0 ),
        .I1(padder_out_1[497]),
        .I2(out[433]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1546]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1290]),
        .O(\out[1229]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1229]_i_3 
       (.I0(\f_permutation_l_/round_in [1393]),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[1229]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[122]_i_1 
       (.I0(\out[1236]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[593] ),
        .I2(\f_permutation_l_/out_reg_n_0_[248] ),
        .I3(\out[1572]_i_3_n_0 ),
        .I4(\out[314]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1230]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1018] ),
        .I1(\out[1416]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[907] ),
        .I3(\out[1230]_i_2_n_0 ),
        .I4(\out[1230]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1230]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1230]_i_2 
       (.I0(\out[1547]_i_16_n_0 ),
        .I1(padder_out_1[498]),
        .I2(out[434]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1547]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1291]),
        .O(\out[1230]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1230]_i_3 
       (.I0(\f_permutation_l_/round_in [1394]),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[1230]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1231]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1019] ),
        .I1(\out[1417]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[908] ),
        .I3(\out[1231]_i_2_n_0 ),
        .I4(\out[1231]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1231]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1231]_i_2 
       (.I0(\out[1548]_i_16_n_0 ),
        .I1(padder_out_1[499]),
        .I2(out[435]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1548]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1292]),
        .O(\out[1231]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1231]_i_3 
       (.I0(\f_permutation_l_/round_in [1395]),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[1231]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1232]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1020] ),
        .I1(\out[1418]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[909] ),
        .I3(\out[1232]_i_2_n_0 ),
        .I4(\out[1232]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1232]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1232]_i_2 
       (.I0(\out[1549]_i_16_n_0 ),
        .I1(padder_out_1[500]),
        .I2(out[436]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1549]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1293]),
        .O(\out[1232]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1232]_i_3 
       (.I0(\f_permutation_l_/round_in [1396]),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[1232]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1233]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1021] ),
        .I1(\out[1419]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[910] ),
        .I3(\out[1233]_i_2_n_0 ),
        .I4(\out[1233]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1233]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1233]_i_2 
       (.I0(\out[1550]_i_16_n_0 ),
        .I1(padder_out_1[501]),
        .I2(out[437]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1550]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1294]),
        .O(\out[1233]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1233]_i_3 
       (.I0(\f_permutation_l_/round_in [1397]),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[1233]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1234]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1022] ),
        .I1(\out[1420]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[911] ),
        .I3(\out[1234]_i_2_n_0 ),
        .I4(\out[1234]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1234]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1234]_i_2 
       (.I0(\out[1551]_i_17_n_0 ),
        .I1(padder_out_1[502]),
        .I2(out[438]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1551]_i_15_n_0 ),
        .I5(\f_permutation_l_/round_in [1295]),
        .O(\out[1234]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1234]_i_3 
       (.I0(\f_permutation_l_/round_in [1398]),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[1234]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1235]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1023] ),
        .I1(\out[1421]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[912] ),
        .I3(\out[1235]_i_2_n_0 ),
        .I4(\out[1235]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1235]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1235]_i_2 
       (.I0(\out[1552]_i_16_n_0 ),
        .I1(padder_out_1[503]),
        .I2(out[439]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1552]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1296]),
        .O(\out[1235]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1235]_i_3 
       (.I0(\f_permutation_l_/round_in [1399]),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[1235]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1236]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[960] ),
        .I1(\out[1422]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[913] ),
        .I3(\out[1236]_i_2_n_0 ),
        .I4(\out[1236]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1236]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1236]_i_2 
       (.I0(\out[1553]_i_16_n_0 ),
        .I1(padder_out_1[488]),
        .I2(out[424]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1553]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1297]),
        .O(\out[1236]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1236]_i_3 
       (.I0(\f_permutation_l_/round_in [1400]),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[1236]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1237]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[961] ),
        .I1(\out[1423]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[914] ),
        .I3(\out[1237]_i_2_n_0 ),
        .I4(\out[1237]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1237]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1237]_i_2 
       (.I0(\out[1554]_i_16_n_0 ),
        .I1(padder_out_1[489]),
        .I2(out[425]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1554]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1298]),
        .O(\out[1237]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1237]_i_3 
       (.I0(\f_permutation_l_/round_in [1401]),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[1237]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1238]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[962] ),
        .I1(\out[1424]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[915] ),
        .I3(\out[1238]_i_2_n_0 ),
        .I4(\out[1238]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1238]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1238]_i_2 
       (.I0(\out[1555]_i_16_n_0 ),
        .I1(padder_out_1[490]),
        .I2(out[426]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1555]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1299]),
        .O(\out[1238]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1238]_i_3 
       (.I0(\f_permutation_l_/round_in [1402]),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[1238]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1239]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[963] ),
        .I1(\out[1425]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[916] ),
        .I3(\out[1239]_i_2_n_0 ),
        .I4(\out[1239]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1239]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1239]_i_2 
       (.I0(\out[1556]_i_16_n_0 ),
        .I1(padder_out_1[491]),
        .I2(out[427]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1556]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1300]),
        .O(\out[1239]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1239]_i_3 
       (.I0(\f_permutation_l_/round_in [1403]),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[1239]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[123]_i_1 
       (.I0(\out[1237]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[594] ),
        .I2(\f_permutation_l_/out_reg_n_0_[249] ),
        .I3(\out[1573]_i_3_n_0 ),
        .I4(\out[315]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1240]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[964] ),
        .I1(\out[1426]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[917] ),
        .I3(\out[1240]_i_2_n_0 ),
        .I4(\out[1240]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1240]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1240]_i_2 
       (.I0(\out[1557]_i_15_n_0 ),
        .I1(padder_out_1[492]),
        .I2(out[428]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1557]_i_13_n_0 ),
        .I5(\f_permutation_l_/round_in [1301]),
        .O(\out[1240]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1240]_i_3 
       (.I0(\f_permutation_l_/round_in [1404]),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[1240]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1241]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[965] ),
        .I1(\out[1427]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[918] ),
        .I3(\out[1241]_i_2_n_0 ),
        .I4(\out[1241]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1241]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1241]_i_2 
       (.I0(\out[1558]_i_14_n_0 ),
        .I1(padder_out_1[302]),
        .I2(out[238]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1493]),
        .I5(\out[1536]_i_14_n_0 ),
        .O(\out[1241]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1241]_i_3 
       (.I0(\f_permutation_l_/round_in [1405]),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[1241]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1242]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[966] ),
        .I1(\out[1428]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[919] ),
        .I3(\out[1242]_i_2_n_0 ),
        .I4(\out[1242]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1242]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1242]_i_2 
       (.I0(\out[1559]_i_15_n_0 ),
        .I1(padder_out_1[303]),
        .I2(out[239]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1537]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1494]),
        .O(\out[1242]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1242]_i_3 
       (.I0(\f_permutation_l_/round_in [1406]),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[1242]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1243]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[967] ),
        .I1(\out[1429]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[920] ),
        .I3(\out[1243]_i_2_n_0 ),
        .I4(\out[1243]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1243]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1243]_i_2 
       (.I0(\out[1560]_i_15_n_0 ),
        .I1(padder_out_1[288]),
        .I2(out[224]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1538]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1495]),
        .O(\out[1243]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1243]_i_3 
       (.I0(\f_permutation_l_/round_in [1407]),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[1243]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1244]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[968] ),
        .I1(\out[1430]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[921] ),
        .I3(\out[1244]_i_2_n_0 ),
        .I4(\out[1244]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1244]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1244]_i_2 
       (.I0(\out[1561]_i_14_n_0 ),
        .I1(padder_out_1[289]),
        .I2(out[225]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1539]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1496]),
        .O(\out[1244]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1244]_i_3 
       (.I0(\f_permutation_l_/round_in [1344]),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[1244]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1245]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[969] ),
        .I1(\out[1431]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[922] ),
        .I3(\out[1245]_i_2_n_0 ),
        .I4(\out[1245]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1245]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1245]_i_2 
       (.I0(\out[1562]_i_15_n_0 ),
        .I1(padder_out_1[290]),
        .I2(out[226]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1540]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1497]),
        .O(\out[1245]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1245]_i_3 
       (.I0(\f_permutation_l_/round_in [1345]),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1409]),
        .I4(\out[1582]_i_7_n_0 ),
        .O(\out[1245]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1246]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[970] ),
        .I1(\out[1432]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[923] ),
        .I3(\out[1246]_i_2_n_0 ),
        .I4(\out[1246]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1246]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1246]_i_2 
       (.I0(\out[1563]_i_14_n_0 ),
        .I1(padder_out_1[291]),
        .I2(out[227]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1541]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1498]),
        .O(\out[1246]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1246]_i_3 
       (.I0(\f_permutation_l_/round_in [1346]),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1410]),
        .I4(\out[1583]_i_7_n_0 ),
        .O(\out[1246]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1247]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[971] ),
        .I1(\out[1433]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[924] ),
        .I3(\out[1247]_i_2_n_0 ),
        .I4(\out[1247]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1247]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1247]_i_2 
       (.I0(\out[1564]_i_15_n_0 ),
        .I1(padder_out_1[292]),
        .I2(out[228]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1542]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1499]),
        .O(\out[1247]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1247]_i_3 
       (.I0(\f_permutation_l_/round_in [1347]),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1411]),
        .I4(\out[1584]_i_7_n_0 ),
        .O(\out[1247]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1248]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[972] ),
        .I1(\out[1434]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[925] ),
        .I3(\out[1248]_i_2_n_0 ),
        .I4(\out[1248]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1248]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1248]_i_2 
       (.I0(\out[1565]_i_15_n_0 ),
        .I1(padder_out_1[293]),
        .I2(out[229]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1543]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1500]),
        .O(\out[1248]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1248]_i_3 
       (.I0(\f_permutation_l_/round_in [1348]),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1412]),
        .I4(\out[1585]_i_7_n_0 ),
        .O(\out[1248]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1249]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[973] ),
        .I1(\out[1435]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[926] ),
        .I3(\out[1249]_i_2_n_0 ),
        .I4(\out[1249]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1249]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1249]_i_2 
       (.I0(\out[1566]_i_14_n_0 ),
        .I1(padder_out_1[294]),
        .I2(out[230]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1544]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1501]),
        .O(\out[1249]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1249]_i_3 
       (.I0(\f_permutation_l_/round_in [1349]),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1413]),
        .I4(\out[1586]_i_7_n_0 ),
        .O(\out[1249]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[124]_i_1 
       (.I0(\out[1238]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[595] ),
        .I2(\f_permutation_l_/out_reg_n_0_[250] ),
        .I3(\out[1574]_i_3_n_0 ),
        .I4(\out[316]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1250]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[974] ),
        .I1(\out[1436]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[927] ),
        .I3(\out[1250]_i_2_n_0 ),
        .I4(\out[1250]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1250]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1250]_i_2 
       (.I0(\out[1567]_i_16_n_0 ),
        .I1(padder_out_1[295]),
        .I2(out[231]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1545]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1502]),
        .O(\out[1250]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1250]_i_3 
       (.I0(\f_permutation_l_/round_in [1350]),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1414]),
        .I4(\out[1587]_i_7_n_0 ),
        .O(\out[1250]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1251]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[975] ),
        .I1(\out[1437]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[928] ),
        .I3(\out[1251]_i_2_n_0 ),
        .I4(\out[1251]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1251]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1251]_i_2 
       (.I0(\out[1568]_i_15_n_0 ),
        .I1(padder_out_1[280]),
        .I2(out[216]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1546]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1503]),
        .O(\out[1251]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1251]_i_3 
       (.I0(\f_permutation_l_/round_in [1351]),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1415]),
        .I4(\out[1588]_i_7_n_0 ),
        .O(\out[1251]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1252]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[976] ),
        .I1(\out[1438]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[929] ),
        .I3(\out[1252]_i_2_n_0 ),
        .I4(\out[1252]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1252]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1252]_i_2 
       (.I0(\out[1569]_i_15_n_0 ),
        .I1(padder_out_1[281]),
        .I2(out[217]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1547]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1504]),
        .O(\out[1252]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1252]_i_3 
       (.I0(\f_permutation_l_/round_in [1352]),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1416]),
        .I4(\out[1589]_i_7_n_0 ),
        .O(\out[1252]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1253]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[977] ),
        .I1(\out[1439]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[930] ),
        .I3(\out[1253]_i_2_n_0 ),
        .I4(\out[1253]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1253]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1253]_i_2 
       (.I0(\out[1570]_i_15_n_0 ),
        .I1(padder_out_1[282]),
        .I2(out[218]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1548]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1505]),
        .O(\out[1253]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1253]_i_3 
       (.I0(\f_permutation_l_/round_in [1353]),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1417]),
        .I4(\out[1590]_i_7_n_0 ),
        .O(\out[1253]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1254]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[978] ),
        .I1(\out[1440]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[931] ),
        .I3(\out[1254]_i_2_n_0 ),
        .I4(\out[1254]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1254]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1254]_i_2 
       (.I0(\out[1571]_i_14_n_0 ),
        .I1(padder_out_1[283]),
        .I2(out[219]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1549]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1506]),
        .O(\out[1254]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1254]_i_3 
       (.I0(\f_permutation_l_/round_in [1354]),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1418]),
        .I4(\out[1591]_i_7_n_0 ),
        .O(\out[1254]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1255]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[979] ),
        .I1(\out[1441]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[932] ),
        .I3(\out[1255]_i_2_n_0 ),
        .I4(\out[1255]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1255]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1255]_i_2 
       (.I0(\out[1572]_i_15_n_0 ),
        .I1(padder_out_1[284]),
        .I2(out[220]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1550]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1507]),
        .O(\out[1255]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1255]_i_3 
       (.I0(\f_permutation_l_/round_in [1355]),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1419]),
        .I4(\out[1592]_i_7_n_0 ),
        .O(\out[1255]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[1256]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[980] ),
        .I1(\out[1442]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[933] ),
        .I3(\out[1256]_i_2_n_0 ),
        .I4(\out[1256]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1256]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1256]_i_2 
       (.I0(\out[1573]_i_15_n_0 ),
        .I1(padder_out_1[285]),
        .I2(out[221]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1551]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1508]),
        .O(\out[1256]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1256]_i_3 
       (.I0(\f_permutation_l_/round_in [1356]),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1420]),
        .I4(\out[1593]_i_7_n_0 ),
        .O(\out[1256]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1257]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[981] ),
        .I1(\out[1443]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[934] ),
        .I3(\out[1257]_i_2_n_0 ),
        .I4(\out[1257]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1257]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1257]_i_2 
       (.I0(\out[1574]_i_15_n_0 ),
        .I1(padder_out_1[286]),
        .I2(out[222]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\out[1552]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1509]),
        .O(\out[1257]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1257]_i_3 
       (.I0(\f_permutation_l_/round_in [1357]),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1421]),
        .I4(\out[1594]_i_7_n_0 ),
        .O(\out[1257]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1258]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[982] ),
        .I1(\out[1444]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[935] ),
        .I3(\out[1258]_i_2_n_0 ),
        .I4(\out[1258]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1258]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1258]_i_2 
       (.I0(\out[1575]_i_15_n_0 ),
        .I1(padder_out_1[287]),
        .I2(out[223]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1553]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1510]),
        .O(\out[1258]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1258]_i_3 
       (.I0(\f_permutation_l_/round_in [1358]),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1422]),
        .I4(\out[1595]_i_7_n_0 ),
        .O(\out[1258]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1259]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[983] ),
        .I1(\out[1445]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[936] ),
        .I3(\out[1259]_i_2_n_0 ),
        .I4(\out[1259]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1259]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1259]_i_2 
       (.I0(\out[1576]_i_15_n_0 ),
        .I1(padder_out_1[272]),
        .I2(out[208]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1554]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1511]),
        .O(\out[1259]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1259]_i_3 
       (.I0(\f_permutation_l_/round_in [1359]),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1423]),
        .I4(\out[1596]_i_7_n_0 ),
        .O(\out[1259]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[125]_i_1 
       (.I0(\out[1239]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[596] ),
        .I2(\f_permutation_l_/out_reg_n_0_[251] ),
        .I3(\out[1575]_i_3_n_0 ),
        .I4(\out[317]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1260]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[984] ),
        .I1(\out[1446]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[937] ),
        .I3(\out[1260]_i_2_n_0 ),
        .I4(\out[1260]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1260]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1260]_i_2 
       (.I0(\out[1577]_i_15_n_0 ),
        .I1(padder_out_1[273]),
        .I2(out[209]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1555]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1512]),
        .O(\out[1260]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1260]_i_3 
       (.I0(\f_permutation_l_/round_in [1360]),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1424]),
        .I4(\out[1597]_i_7_n_0 ),
        .O(\out[1260]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1261]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[985] ),
        .I1(\out[1447]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[938] ),
        .I3(\out[1261]_i_2_n_0 ),
        .I4(\out[1261]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1261]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1261]_i_2 
       (.I0(\out[1578]_i_14_n_0 ),
        .I1(padder_out_1[274]),
        .I2(out[210]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1556]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1513]),
        .O(\out[1261]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1261]_i_3 
       (.I0(\f_permutation_l_/round_in [1361]),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1425]),
        .I4(\out[1598]_i_7_n_0 ),
        .O(\out[1261]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1262]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[986] ),
        .I1(\out[1448]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[939] ),
        .I3(\out[1262]_i_2_n_0 ),
        .I4(\out[1262]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1262]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1262]_i_2 
       (.I0(\out[1579]_i_15_n_0 ),
        .I1(padder_out_1[275]),
        .I2(out[211]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1557]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1514]),
        .O(\out[1262]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1262]_i_3 
       (.I0(\f_permutation_l_/round_in [1362]),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\out[1599]_i_7_n_0 ),
        .I4(\f_permutation_l_/round_in [1426]),
        .O(\out[1262]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1263]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[987] ),
        .I1(\out[1449]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[940] ),
        .I3(\out[1263]_i_2_n_0 ),
        .I4(\out[1263]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1263]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1263]_i_2 
       (.I0(\out[1580]_i_14_n_0 ),
        .I1(padder_out_1[276]),
        .I2(out[212]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1558]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1515]),
        .O(\out[1263]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1263]_i_3 
       (.I0(\f_permutation_l_/round_in [1363]),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\out[1554]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1298]),
        .O(\out[1263]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1264]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[988] ),
        .I1(\out[1450]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[941] ),
        .I3(\out[1264]_i_2_n_0 ),
        .I4(\out[1264]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1264]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1264]_i_2 
       (.I0(\out[1581]_i_14_n_0 ),
        .I1(padder_out_1[277]),
        .I2(out[213]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1559]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1516]),
        .O(\out[1264]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1264]_i_3 
       (.I0(\f_permutation_l_/round_in [1364]),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\out[1555]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1299]),
        .O(\out[1264]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1265]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[989] ),
        .I1(\out[1451]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[942] ),
        .I3(\out[1265]_i_2_n_0 ),
        .I4(\out[1265]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1265]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1265]_i_2 
       (.I0(\out[1582]_i_14_n_0 ),
        .I1(padder_out_1[278]),
        .I2(out[214]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1560]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1517]),
        .O(\out[1265]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1265]_i_3 
       (.I0(\f_permutation_l_/round_in [1365]),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\out[1556]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1300]),
        .O(\out[1265]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1266]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[990] ),
        .I1(\out[1452]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[943] ),
        .I3(\out[1266]_i_2_n_0 ),
        .I4(\out[1266]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1266]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1266]_i_2 
       (.I0(\out[1583]_i_14_n_0 ),
        .I1(padder_out_1[279]),
        .I2(out[215]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1561]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1518]),
        .O(\out[1266]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1266]_i_3 
       (.I0(\f_permutation_l_/round_in [1366]),
        .I1(\f_permutation_l_/round_in [1430]),
        .I2(\out[1539]_i_9_n_0 ),
        .I3(\out[1557]_i_13_n_0 ),
        .I4(\f_permutation_l_/round_in [1301]),
        .O(\out[1266]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1267]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[991] ),
        .I1(\out[1453]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[944] ),
        .I3(\out[1267]_i_2_n_0 ),
        .I4(\out[1267]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1267]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1267]_i_2 
       (.I0(\out[1584]_i_14_n_0 ),
        .I1(padder_out_1[264]),
        .I2(out[200]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1562]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1519]),
        .O(\out[1267]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1267]_i_3 
       (.I0(\f_permutation_l_/round_in [1367]),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[1267]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1268]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[992] ),
        .I1(\out[1454]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[945] ),
        .I3(\out[1268]_i_2_n_0 ),
        .I4(\out[1268]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1268]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1268]_i_2 
       (.I0(\out[1585]_i_14_n_0 ),
        .I1(padder_out_1[265]),
        .I2(out[201]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1563]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1520]),
        .O(\out[1268]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1268]_i_3 
       (.I0(\f_permutation_l_/round_in [1368]),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[1268]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1269]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[993] ),
        .I1(\out[1455]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[946] ),
        .I3(\out[1269]_i_2_n_0 ),
        .I4(\out[1269]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1269]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1269]_i_2 
       (.I0(\out[1586]_i_14_n_0 ),
        .I1(padder_out_1[266]),
        .I2(out[202]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1564]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1521]),
        .O(\out[1269]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1269]_i_3 
       (.I0(\f_permutation_l_/round_in [1369]),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[1269]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[126]_i_1 
       (.I0(\out[1240]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[597] ),
        .I2(\f_permutation_l_/out_reg_n_0_[252] ),
        .I3(\out[1576]_i_3_n_0 ),
        .I4(\out[318]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1270]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[994] ),
        .I1(\out[1456]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[947] ),
        .I3(\out[1270]_i_2_n_0 ),
        .I4(\out[1270]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1270]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1270]_i_2 
       (.I0(\out[1587]_i_13_n_0 ),
        .I1(padder_out_1[267]),
        .I2(out[203]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1565]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1522]),
        .O(\out[1270]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1270]_i_3 
       (.I0(\f_permutation_l_/round_in [1370]),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[1270]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1271]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[995] ),
        .I1(\out[1457]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[948] ),
        .I3(\out[1271]_i_2_n_0 ),
        .I4(\out[1271]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1271]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1271]_i_2 
       (.I0(\out[1588]_i_14_n_0 ),
        .I1(padder_out_1[268]),
        .I2(out[204]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1566]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1523]),
        .O(\out[1271]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1271]_i_3 
       (.I0(\f_permutation_l_/round_in [1371]),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[1271]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1272]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[996] ),
        .I1(\out[1458]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[949] ),
        .I3(\out[1272]_i_2_n_0 ),
        .I4(\out[1272]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1272]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1272]_i_2 
       (.I0(\out[1589]_i_14_n_0 ),
        .I1(padder_out_1[269]),
        .I2(out[205]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1567]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1524]),
        .O(\out[1272]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1272]_i_3 
       (.I0(\f_permutation_l_/round_in [1372]),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[1272]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1273]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[997] ),
        .I1(\out[1459]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[950] ),
        .I3(\out[1273]_i_2_n_0 ),
        .I4(\out[1273]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1273]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1273]_i_2 
       (.I0(\out[1590]_i_14_n_0 ),
        .I1(padder_out_1[270]),
        .I2(out[206]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1568]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1525]),
        .O(\out[1273]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1273]_i_3 
       (.I0(\f_permutation_l_/round_in [1373]),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[1273]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1274]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[998] ),
        .I1(\out[1460]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[951] ),
        .I3(\out[1274]_i_2_n_0 ),
        .I4(\out[1274]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1274]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1274]_i_2 
       (.I0(\out[1591]_i_14_n_0 ),
        .I1(padder_out_1[271]),
        .I2(out[207]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1569]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1526]),
        .O(\out[1274]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1274]_i_3 
       (.I0(\f_permutation_l_/round_in [1374]),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[1274]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1275]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[999] ),
        .I1(\out[1461]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[952] ),
        .I3(\out[1275]_i_2_n_0 ),
        .I4(\out[1275]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1275]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1275]_i_2 
       (.I0(\out[1592]_i_14_n_0 ),
        .I1(padder_out_1[256]),
        .I2(out[192]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1570]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1527]),
        .O(\out[1275]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1275]_i_3 
       (.I0(\f_permutation_l_/round_in [1375]),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[1275]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1276]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1000] ),
        .I1(\out[1462]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[953] ),
        .I3(\out[1276]_i_2_n_0 ),
        .I4(\out[1276]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1276]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1276]_i_2 
       (.I0(\out[1593]_i_14_n_0 ),
        .I1(padder_out_1[257]),
        .I2(out[193]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1571]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1528]),
        .O(\out[1276]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1276]_i_3 
       (.I0(\f_permutation_l_/round_in [1376]),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[1276]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1277]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1001] ),
        .I1(\out[1463]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[954] ),
        .I3(\out[1277]_i_2_n_0 ),
        .I4(\out[1277]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1277]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1277]_i_2 
       (.I0(\out[1594]_i_14_n_0 ),
        .I1(padder_out_1[258]),
        .I2(out[194]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1572]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1529]),
        .O(\out[1277]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1277]_i_3 
       (.I0(\f_permutation_l_/round_in [1377]),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[1277]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1278]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1002] ),
        .I1(\out[1464]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[955] ),
        .I3(\out[1278]_i_2_n_0 ),
        .I4(\out[1278]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1278]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1278]_i_2 
       (.I0(\out[1595]_i_14_n_0 ),
        .I1(padder_out_1[259]),
        .I2(out[195]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1573]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1530]),
        .O(\out[1278]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1278]_i_3 
       (.I0(\f_permutation_l_/round_in [1378]),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[1278]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1279]_i_1 
       (.I0(\f_permutation_l_/out_reg_n_0_[1003] ),
        .I1(\out[1465]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[956] ),
        .I3(\out[1279]_i_2_n_0 ),
        .I4(\out[1279]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1279]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1279]_i_2 
       (.I0(\out[1596]_i_14_n_0 ),
        .I1(padder_out_1[260]),
        .I2(out[196]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\out[1574]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1531]),
        .O(\out[1279]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1279]_i_3 
       (.I0(\f_permutation_l_/round_in [1379]),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[1279]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[127]_i_1 
       (.I0(\out[1241]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[598] ),
        .I2(\f_permutation_l_/out_reg_n_0_[253] ),
        .I3(\out[1577]_i_3_n_0 ),
        .I4(\out[319]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1280]_i_1 
       (.I0(\out[1408]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[50] ),
        .I2(\out[1536]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1172]),
        .I4(\out[1280]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1280]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1280]_i_2 
       (.I0(padder_out_1[172]),
        .I1(out[108]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1172]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1280]_i_3 
       (.I0(\out[1536]_i_10_n_0 ),
        .I1(padder_out_1[556]),
        .I2(out[492]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1536]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1427]),
        .O(\out[1280]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1281]_i_1 
       (.I0(\out[1409]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[51] ),
        .I2(\out[1537]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1173]),
        .I4(\out[1281]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1281]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1281]_i_2 
       (.I0(padder_out_1[173]),
        .I1(out[109]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1173]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1281]_i_3 
       (.I0(\out[1537]_i_9_n_0 ),
        .I1(padder_out_1[557]),
        .I2(out[493]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1537]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1428]),
        .O(\out[1281]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1282]_i_1 
       (.I0(\out[1410]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[52] ),
        .I2(\out[1538]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1174]),
        .I4(\out[1538]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1282]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1283]_i_1 
       (.I0(\out[1411]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[53] ),
        .I2(\out[1347]_i_2_n_0 ),
        .I3(\f_permutation_l_/round_in [1175]),
        .I4(\out[1539]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1283]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1284]_i_1 
       (.I0(\out[1412]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[54] ),
        .I2(\out[1540]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1176]),
        .I4(\out[1540]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1284]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1285]_i_1 
       (.I0(\out[1413]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[55] ),
        .I2(\out[1541]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1177]),
        .I4(\out[1541]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1285]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1286]_i_1 
       (.I0(\out[1414]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[56] ),
        .I2(\out[1542]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1178]),
        .I4(\out[1542]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1286]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1287]_i_1 
       (.I0(\out[1415]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[57] ),
        .I2(\out[1543]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1179]),
        .I4(\out[1287]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1287]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1287]_i_2 
       (.I0(padder_out_1[163]),
        .I1(out[99]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1179]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1287]_i_3 
       (.I0(\out[1543]_i_10_n_0 ),
        .I1(padder_out_1[547]),
        .I2(out[483]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1543]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1434]),
        .O(\out[1287]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1288]_i_1 
       (.I0(\out[1416]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[58] ),
        .I2(\out[1544]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1180]),
        .I4(\out[1544]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1288]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1289]_i_1 
       (.I0(\out[1417]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[59] ),
        .I2(\out[1545]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1181]),
        .I4(\out[1545]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1289]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[128]_i_1 
       (.I0(\out[1447]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[665] ),
        .I2(\out[128]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[254] ),
        .I4(\out[1578]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [128]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[128]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[599] ),
        .I1(\f_permutation_l_/round_in [1494]),
        .I2(\out[1537]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[128]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1290]_i_1 
       (.I0(\out[1418]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[60] ),
        .I2(\out[1546]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1182]),
        .I4(\out[1546]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1290]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1291]_i_1 
       (.I0(\out[1419]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[61] ),
        .I2(\out[1547]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1183]),
        .I4(\out[1547]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1291]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1292]_i_1 
       (.I0(\out[1420]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[62] ),
        .I2(\out[1548]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1184]),
        .I4(\out[1548]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1292]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1293]_i_1 
       (.I0(\out[1421]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[63] ),
        .I2(\out[1549]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1185]),
        .I4(\out[1549]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1293]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1294]_i_1 
       (.I0(\out[1422]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_ ),
        .I2(\out[1550]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1186]),
        .I4(\out[1550]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1294]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1295]_i_1 
       (.I0(\out[1423]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[1] ),
        .I2(\out[1551]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1187]),
        .I4(\out[1295]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1295]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1295]_i_2 
       (.I0(padder_out_1[155]),
        .I1(out[91]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1187]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1295]_i_3 
       (.I0(\out[1551]_i_9_n_0 ),
        .I1(padder_out_1[539]),
        .I2(out[475]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1551]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1442]),
        .O(\out[1295]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1296]_i_1 
       (.I0(\out[1424]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[2] ),
        .I2(\out[1552]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1188]),
        .I4(\out[1552]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1296]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1297]_i_1 
       (.I0(\out[1425]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[3] ),
        .I2(\out[1553]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1189]),
        .I4(\out[1553]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1297]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1298]_i_1 
       (.I0(\out[1426]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[4] ),
        .I2(\out[1554]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1190]),
        .I4(\out[1554]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1298]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1299]_i_1 
       (.I0(\out[1427]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[5] ),
        .I2(\out[1555]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1191]),
        .I4(\out[1555]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1299]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[129]_i_1 
       (.I0(\out[1448]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[666] ),
        .I2(\out[129]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[255] ),
        .I4(\out[1579]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [129]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[129]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[600] ),
        .I1(\f_permutation_l_/round_in [1495]),
        .I2(\out[1538]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[129]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[12]_i_1 
       (.I0(\out[1590]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[202] ),
        .I2(\out[268]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1045]),
        .I4(\out[1514]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1300]_i_1 
       (.I0(\out[1428]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[6] ),
        .I2(\out[1556]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1192]),
        .I4(\out[1556]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1300]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1301]_i_1 
       (.I0(\out[1429]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[7] ),
        .I2(\out[1557]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1193]),
        .I4(\out[1557]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1301]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1302]_i_1 
       (.I0(\out[1430]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[8] ),
        .I2(\out[1558]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1194]),
        .I4(\out[1558]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1302]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1303]_i_1 
       (.I0(\out[1431]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[9] ),
        .I2(\out[1559]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1195]),
        .I4(\out[1559]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1303]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1304]_i_1 
       (.I0(\out[1432]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[10] ),
        .I2(\out[1560]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1196]),
        .I4(\out[1560]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1304]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1305]_i_1 
       (.I0(\out[1433]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[11] ),
        .I2(\out[1561]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1197]),
        .I4(\out[1561]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1305]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1306]_i_1 
       (.I0(\out[1434]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[12] ),
        .I2(\out[1562]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1198]),
        .I4(\out[1562]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1306]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1307]_i_1 
       (.I0(\out[1435]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[13] ),
        .I2(\out[1563]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1199]),
        .I4(\out[1563]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1307]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1308]_i_1 
       (.I0(\out[1436]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[14] ),
        .I2(\out[1564]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1200]),
        .I4(\out[1564]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1308]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1309]_i_1 
       (.I0(\out[1437]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[15] ),
        .I2(\out[1565]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1201]),
        .I4(\out[1565]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1309]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[130]_i_1 
       (.I0(\out[1449]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[667] ),
        .I2(\out[130]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[192] ),
        .I4(\out[1580]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [130]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[130]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[601] ),
        .I1(\f_permutation_l_/round_in [1496]),
        .I2(\out[1539]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[130]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1310]_i_1 
       (.I0(\out[1438]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[16] ),
        .I2(\out[1566]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1202]),
        .I4(\out[1566]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1310]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1311]_i_1 
       (.I0(\out[1439]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[17] ),
        .I2(\out[1567]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1203]),
        .I4(\out[1311]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1311]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1311]_i_2 
       (.I0(padder_out_1[139]),
        .I1(out[75]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1203]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1311]_i_3 
       (.I0(\out[1567]_i_9_n_0 ),
        .I1(padder_out_1[523]),
        .I2(out[459]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1567]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1458]),
        .O(\out[1311]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1312]_i_1 
       (.I0(\out[1440]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[18] ),
        .I2(\out[1568]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1204]),
        .I4(\out[1568]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1312]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1313]_i_1 
       (.I0(\out[1441]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[19] ),
        .I2(\out[1569]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1205]),
        .I4(\out[1569]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1313]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1314]_i_1 
       (.I0(\out[1442]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[20] ),
        .I2(\out[1570]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1206]),
        .I4(\out[1570]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1314]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1315]_i_1 
       (.I0(\out[1443]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[21] ),
        .I2(\out[1571]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1207]),
        .I4(\out[1571]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1315]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1316]_i_1 
       (.I0(\out[1444]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[22] ),
        .I2(\out[1572]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1208]),
        .I4(\out[1572]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1316]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1317]_i_1 
       (.I0(\out[1445]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[23] ),
        .I2(\out[1573]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1209]),
        .I4(\out[1573]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1317]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1318]_i_1 
       (.I0(\out[1446]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[24] ),
        .I2(\out[1574]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1210]),
        .I4(\out[1574]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1318]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1319]_i_1 
       (.I0(\out[1447]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[25] ),
        .I2(\out[1575]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1211]),
        .I4(\out[1575]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1319]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[131]_i_1 
       (.I0(\out[1450]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[668] ),
        .I2(\out[131]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[193] ),
        .I4(\out[1581]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [131]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[131]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[602] ),
        .I1(\f_permutation_l_/round_in [1497]),
        .I2(\out[1540]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[131]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1320]_i_1 
       (.I0(\out[1448]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[26] ),
        .I2(\out[1576]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1212]),
        .I4(\out[1576]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1320]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1321]_i_1 
       (.I0(\out[1449]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[27] ),
        .I2(\out[1577]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1213]),
        .I4(\out[1577]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1321]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1322]_i_1 
       (.I0(\out[1450]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[28] ),
        .I2(\out[1578]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1214]),
        .I4(\out[1578]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1322]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1323]_i_1 
       (.I0(\out[1451]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[29] ),
        .I2(\out[1579]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1215]),
        .I4(\out[1579]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1323]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1324]_i_1 
       (.I0(\out[1452]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[30] ),
        .I2(\out[1580]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1152]),
        .I4(\out[1580]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1324]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1325]_i_1 
       (.I0(\out[1453]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[31] ),
        .I2(\out[1581]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1153]),
        .I4(\out[1581]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1325]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1326]_i_1 
       (.I0(\out[1454]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[32] ),
        .I2(\out[1582]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1154]),
        .I4(\out[1582]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1326]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1327]_i_1 
       (.I0(\out[1455]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[33] ),
        .I2(\out[1583]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1155]),
        .I4(\out[1583]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1327]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1328]_i_1 
       (.I0(\out[1456]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[34] ),
        .I2(\out[1584]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1156]),
        .I4(\out[1584]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1328]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1329]_i_1 
       (.I0(\out[1457]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[35] ),
        .I2(\out[1585]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1157]),
        .I4(\out[1585]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1329]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[132]_i_1 
       (.I0(\out[1451]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[669] ),
        .I2(\out[132]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[194] ),
        .I4(\out[1582]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [132]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[132]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[603] ),
        .I1(\f_permutation_l_/round_in [1498]),
        .I2(\out[1541]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[132]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1330]_i_1 
       (.I0(\out[1458]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[36] ),
        .I2(\out[1586]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1158]),
        .I4(\out[1586]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1330]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1331]_i_1 
       (.I0(\out[1459]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[37] ),
        .I2(\out[1587]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1159]),
        .I4(\out[1587]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1331]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1332]_i_1 
       (.I0(\out[1460]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[38] ),
        .I2(\out[1588]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1160]),
        .I4(\out[1588]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1332]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1333]_i_1 
       (.I0(\out[1461]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[39] ),
        .I2(\out[1589]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1161]),
        .I4(\out[1589]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1333]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1334]_i_1 
       (.I0(\out[1462]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[40] ),
        .I2(\out[1590]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1162]),
        .I4(\out[1590]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1334]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1335]_i_1 
       (.I0(\out[1463]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[41] ),
        .I2(\out[1591]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1163]),
        .I4(\out[1591]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1335]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1336]_i_1 
       (.I0(\out[1464]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[42] ),
        .I2(\out[1592]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1164]),
        .I4(\out[1592]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1336]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1337]_i_1 
       (.I0(\out[1465]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[43] ),
        .I2(\out[1593]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1165]),
        .I4(\out[1593]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1337]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1338]_i_1 
       (.I0(\out[1466]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[44] ),
        .I2(\out[1594]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1166]),
        .I4(\out[1594]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1338]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1339]_i_1 
       (.I0(\out[1467]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[45] ),
        .I2(\out[1595]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1167]),
        .I4(\out[1595]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1339]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[133]_i_1 
       (.I0(\out[1452]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[670] ),
        .I2(\out[133]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[195] ),
        .I4(\out[1583]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [133]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[133]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[604] ),
        .I1(\f_permutation_l_/round_in [1499]),
        .I2(\out[1542]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[133]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1340]_i_1 
       (.I0(\out[1468]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[46] ),
        .I2(\out[1596]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1168]),
        .I4(\out[1596]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1340]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1341]_i_1 
       (.I0(\out[1469]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[47] ),
        .I2(\out[1597]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1169]),
        .I4(\out[1597]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1341]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1342]_i_1 
       (.I0(\out[1470]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[48] ),
        .I2(\out[1598]_i_5_n_0 ),
        .I3(\f_permutation_l_/round_in [1170]),
        .I4(\out[1598]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1342]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1343]_i_1 
       (.I0(\out[1471]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[49] ),
        .I2(\out[1599]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1171]),
        .I4(\out[1343]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1343]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1343]_i_2 
       (.I0(padder_out_1[171]),
        .I1(out[107]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1171]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1343]_i_3 
       (.I0(\out[1599]_i_8_n_0 ),
        .I1(padder_out_1[555]),
        .I2(out[491]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1599]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1426]),
        .O(\out[1343]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1344]_i_1 
       (.I0(\out[1472]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[427] ),
        .I2(\f_permutation_l_/out_reg_n_0_[50] ),
        .I3(\out[1408]_i_3_n_0 ),
        .I4(\out[1536]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1344]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1345]_i_1 
       (.I0(\out[1473]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[428] ),
        .I2(\f_permutation_l_/out_reg_n_0_[51] ),
        .I3(\out[1409]_i_3_n_0 ),
        .I4(\out[1537]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1345]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1346]_i_1 
       (.I0(\out[1474]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[429] ),
        .I2(\f_permutation_l_/out_reg_n_0_[52] ),
        .I3(\out[1410]_i_3_n_0 ),
        .I4(\out[1538]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1346]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1347]_i_1 
       (.I0(\out[1475]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[430] ),
        .I2(\f_permutation_l_/out_reg_n_0_[53] ),
        .I3(\out[1411]_i_2_n_0 ),
        .I4(\out[1347]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1347]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1347]_i_2 
       (.I0(\f_permutation_l_/round_in [1539]),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[1347]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1347]_i_3 
       (.I0(padder_out_1[506]),
        .I1(out[442]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1474]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1348]_i_1 
       (.I0(\out[1476]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[431] ),
        .I2(\f_permutation_l_/out_reg_n_0_[54] ),
        .I3(\out[1412]_i_3_n_0 ),
        .I4(\out[1540]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1348]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1349]_i_1 
       (.I0(\out[1477]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[432] ),
        .I2(\f_permutation_l_/out_reg_n_0_[55] ),
        .I3(\out[1413]_i_3_n_0 ),
        .I4(\out[1541]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1349]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[134]_i_1 
       (.I0(\out[1453]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[671] ),
        .I2(\out[134]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[196] ),
        .I4(\out[1584]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [134]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[134]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[605] ),
        .I1(\f_permutation_l_/round_in [1500]),
        .I2(\out[1543]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[134]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1350]_i_1 
       (.I0(\out[1478]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[433] ),
        .I2(\f_permutation_l_/out_reg_n_0_[56] ),
        .I3(\out[1414]_i_3_n_0 ),
        .I4(\out[1542]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1350]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1351]_i_1 
       (.I0(\out[1479]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[434] ),
        .I2(\f_permutation_l_/out_reg_n_0_[57] ),
        .I3(\out[1415]_i_3_n_0 ),
        .I4(\out[1543]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1351]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1352]_i_1 
       (.I0(\out[1480]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[435] ),
        .I2(\f_permutation_l_/out_reg_n_0_[58] ),
        .I3(\out[1416]_i_3_n_0 ),
        .I4(\out[1544]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1352]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1353]_i_1 
       (.I0(\out[1481]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[436] ),
        .I2(\f_permutation_l_/out_reg_n_0_[59] ),
        .I3(\out[1417]_i_3_n_0 ),
        .I4(\out[1545]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1353]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1354]_i_1 
       (.I0(\out[1482]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[437] ),
        .I2(\f_permutation_l_/out_reg_n_0_[60] ),
        .I3(\out[1418]_i_3_n_0 ),
        .I4(\out[1546]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1354]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1355]_i_1 
       (.I0(\out[1483]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[438] ),
        .I2(\f_permutation_l_/out_reg_n_0_[61] ),
        .I3(\out[1419]_i_3_n_0 ),
        .I4(\out[1547]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1355]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1356]_i_1 
       (.I0(\out[1484]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[439] ),
        .I2(\f_permutation_l_/out_reg_n_0_[62] ),
        .I3(\out[1420]_i_3_n_0 ),
        .I4(\out[1548]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1356]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1357]_i_1 
       (.I0(\out[1485]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[440] ),
        .I2(\f_permutation_l_/out_reg_n_0_[63] ),
        .I3(\out[1421]_i_3_n_0 ),
        .I4(\out[1549]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1357]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1358]_i_1 
       (.I0(\out[1486]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[441] ),
        .I2(\f_permutation_l_/out_reg_n_0_ ),
        .I3(\out[1422]_i_3_n_0 ),
        .I4(\out[1550]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1358]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1359]_i_1 
       (.I0(\out[1487]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[442] ),
        .I2(\f_permutation_l_/out_reg_n_0_[1] ),
        .I3(\out[1423]_i_3_n_0 ),
        .I4(\out[1551]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1359]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[135]_i_1 
       (.I0(\out[1454]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[672] ),
        .I2(\out[135]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[197] ),
        .I4(\out[1585]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [135]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[135]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[606] ),
        .I1(\f_permutation_l_/round_in [1501]),
        .I2(\out[1544]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[135]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1360]_i_1 
       (.I0(\out[1488]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[443] ),
        .I2(\f_permutation_l_/out_reg_n_0_[2] ),
        .I3(\out[1424]_i_3_n_0 ),
        .I4(\out[1552]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1360]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1361]_i_1 
       (.I0(\out[1489]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[444] ),
        .I2(\f_permutation_l_/out_reg_n_0_[3] ),
        .I3(\out[1425]_i_3_n_0 ),
        .I4(\out[1553]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1361]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1362]_i_1 
       (.I0(\out[1490]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[445] ),
        .I2(\f_permutation_l_/out_reg_n_0_[4] ),
        .I3(\out[1426]_i_3_n_0 ),
        .I4(\out[1554]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1362]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1363]_i_1 
       (.I0(\out[1491]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[446] ),
        .I2(\f_permutation_l_/out_reg_n_0_[5] ),
        .I3(\out[1427]_i_3_n_0 ),
        .I4(\out[1555]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1363]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1364]_i_1 
       (.I0(\out[1492]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[447] ),
        .I2(\f_permutation_l_/out_reg_n_0_[6] ),
        .I3(\out[1428]_i_3_n_0 ),
        .I4(\out[1556]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1364]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1365]_i_1 
       (.I0(\out[1493]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[384] ),
        .I2(\f_permutation_l_/out_reg_n_0_[7] ),
        .I3(\out[1429]_i_3_n_0 ),
        .I4(\out[1557]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1365]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1366]_i_1 
       (.I0(\out[1494]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[385] ),
        .I2(\f_permutation_l_/out_reg_n_0_[8] ),
        .I3(\out[1430]_i_3_n_0 ),
        .I4(\out[1558]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1366]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1367]_i_1 
       (.I0(\out[1495]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[386] ),
        .I2(\f_permutation_l_/out_reg_n_0_[9] ),
        .I3(\out[1431]_i_3_n_0 ),
        .I4(\out[1559]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1367]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1368]_i_1 
       (.I0(\out[1496]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[387] ),
        .I2(\f_permutation_l_/out_reg_n_0_[10] ),
        .I3(\out[1432]_i_3_n_0 ),
        .I4(\out[1560]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1368]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1369]_i_1 
       (.I0(\out[1497]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[388] ),
        .I2(\f_permutation_l_/out_reg_n_0_[11] ),
        .I3(\out[1433]_i_3_n_0 ),
        .I4(\out[1561]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1369]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[136]_i_1 
       (.I0(\out[1455]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[673] ),
        .I2(\out[136]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[198] ),
        .I4(\out[1586]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [136]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[136]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[607] ),
        .I1(\f_permutation_l_/round_in [1502]),
        .I2(\out[1545]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[136]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1370]_i_1 
       (.I0(\out[1498]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[389] ),
        .I2(\f_permutation_l_/out_reg_n_0_[12] ),
        .I3(\out[1434]_i_3_n_0 ),
        .I4(\out[1562]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1370]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1371]_i_1 
       (.I0(\out[1499]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[390] ),
        .I2(\f_permutation_l_/out_reg_n_0_[13] ),
        .I3(\out[1435]_i_3_n_0 ),
        .I4(\out[1563]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1371]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1372]_i_1 
       (.I0(\out[1500]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[391] ),
        .I2(\f_permutation_l_/out_reg_n_0_[14] ),
        .I3(\out[1436]_i_3_n_0 ),
        .I4(\out[1564]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1372]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1373]_i_1 
       (.I0(\out[1501]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[392] ),
        .I2(\f_permutation_l_/out_reg_n_0_[15] ),
        .I3(\out[1437]_i_3_n_0 ),
        .I4(\out[1565]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1373]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1374]_i_1 
       (.I0(\out[1502]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[393] ),
        .I2(\f_permutation_l_/out_reg_n_0_[16] ),
        .I3(\out[1438]_i_3_n_0 ),
        .I4(\out[1566]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1374]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1375]_i_1 
       (.I0(\out[1503]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[394] ),
        .I2(\f_permutation_l_/out_reg_n_0_[17] ),
        .I3(\out[1439]_i_3_n_0 ),
        .I4(\out[1567]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1375]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1376]_i_1 
       (.I0(\out[1504]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[395] ),
        .I2(\f_permutation_l_/out_reg_n_0_[18] ),
        .I3(\out[1440]_i_3_n_0 ),
        .I4(\out[1568]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1376]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1377]_i_1 
       (.I0(\out[1505]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[396] ),
        .I2(\f_permutation_l_/out_reg_n_0_[19] ),
        .I3(\out[1441]_i_3_n_0 ),
        .I4(\out[1569]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1377]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[1378]_i_1 
       (.I0(\out[1506]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[397] ),
        .I2(\f_permutation_l_/out_reg_n_0_[20] ),
        .I3(\out[1442]_i_3_n_0 ),
        .I4(\out[1570]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1378]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1379]_i_1 
       (.I0(\out[1507]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[398] ),
        .I2(\f_permutation_l_/out_reg_n_0_[21] ),
        .I3(\out[1443]_i_3_n_0 ),
        .I4(\out[1571]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1379]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[137]_i_1 
       (.I0(\out[1456]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[674] ),
        .I2(\out[137]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[199] ),
        .I4(\out[1587]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [137]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[137]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[608] ),
        .I1(\f_permutation_l_/round_in [1503]),
        .I2(\out[1546]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[137]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1380]_i_1 
       (.I0(\out[1508]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[399] ),
        .I2(\f_permutation_l_/out_reg_n_0_[22] ),
        .I3(\out[1444]_i_3_n_0 ),
        .I4(\out[1572]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1380]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1381]_i_1 
       (.I0(\out[1509]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[400] ),
        .I2(\f_permutation_l_/out_reg_n_0_[23] ),
        .I3(\out[1445]_i_3_n_0 ),
        .I4(\out[1573]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1381]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1382]_i_1 
       (.I0(\out[1510]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[401] ),
        .I2(\f_permutation_l_/out_reg_n_0_[24] ),
        .I3(\out[1446]_i_3_n_0 ),
        .I4(\out[1574]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1382]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1383]_i_1 
       (.I0(\out[1511]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[402] ),
        .I2(\f_permutation_l_/out_reg_n_0_[25] ),
        .I3(\out[1447]_i_3_n_0 ),
        .I4(\out[1575]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1383]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1384]_i_1 
       (.I0(\out[1512]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[403] ),
        .I2(\f_permutation_l_/out_reg_n_0_[26] ),
        .I3(\out[1448]_i_3_n_0 ),
        .I4(\out[1576]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1384]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1385]_i_1 
       (.I0(\out[1513]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[404] ),
        .I2(\f_permutation_l_/out_reg_n_0_[27] ),
        .I3(\out[1449]_i_3_n_0 ),
        .I4(\out[1577]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1385]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1386]_i_1 
       (.I0(\out[1514]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[405] ),
        .I2(\f_permutation_l_/out_reg_n_0_[28] ),
        .I3(\out[1450]_i_3_n_0 ),
        .I4(\out[1578]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1386]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[1387]_i_1 
       (.I0(\out[1515]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[406] ),
        .I2(\f_permutation_l_/out_reg_n_0_[29] ),
        .I3(\out[1451]_i_3_n_0 ),
        .I4(\out[1579]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1387]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1388]_i_1 
       (.I0(\out[1516]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[407] ),
        .I2(\f_permutation_l_/out_reg_n_0_[30] ),
        .I3(\out[1452]_i_3_n_0 ),
        .I4(\out[1580]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1388]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1389]_i_1 
       (.I0(\out[1517]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[408] ),
        .I2(\f_permutation_l_/out_reg_n_0_[31] ),
        .I3(\out[1453]_i_3_n_0 ),
        .I4(\out[1581]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1389]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[138]_i_1 
       (.I0(\out[1457]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[675] ),
        .I2(\out[138]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[200] ),
        .I4(\out[1588]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [138]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[138]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[609] ),
        .I1(\f_permutation_l_/round_in [1504]),
        .I2(\out[1547]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[138]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1390]_i_1 
       (.I0(\out[1518]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[409] ),
        .I2(\f_permutation_l_/out_reg_n_0_[32] ),
        .I3(\out[1454]_i_3_n_0 ),
        .I4(\out[1582]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1390]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1391]_i_1 
       (.I0(\out[1519]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[410] ),
        .I2(\f_permutation_l_/out_reg_n_0_[33] ),
        .I3(\out[1455]_i_3_n_0 ),
        .I4(\out[1583]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1391]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1392]_i_1 
       (.I0(\out[1520]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[411] ),
        .I2(\f_permutation_l_/out_reg_n_0_[34] ),
        .I3(\out[1456]_i_3_n_0 ),
        .I4(\out[1584]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1392]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1393]_i_1 
       (.I0(\out[1521]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[412] ),
        .I2(\f_permutation_l_/out_reg_n_0_[35] ),
        .I3(\out[1457]_i_3_n_0 ),
        .I4(\out[1585]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1393]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1394]_i_1 
       (.I0(\out[1522]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[413] ),
        .I2(\f_permutation_l_/out_reg_n_0_[36] ),
        .I3(\out[1458]_i_3_n_0 ),
        .I4(\out[1586]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1394]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1395]_i_1 
       (.I0(\out[1523]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[414] ),
        .I2(\f_permutation_l_/out_reg_n_0_[37] ),
        .I3(\out[1459]_i_3_n_0 ),
        .I4(\out[1587]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1395]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1396]_i_1 
       (.I0(\out[1524]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[415] ),
        .I2(\f_permutation_l_/out_reg_n_0_[38] ),
        .I3(\out[1460]_i_3_n_0 ),
        .I4(\out[1588]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1396]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1397]_i_1 
       (.I0(\out[1525]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[416] ),
        .I2(\f_permutation_l_/out_reg_n_0_[39] ),
        .I3(\out[1461]_i_3_n_0 ),
        .I4(\out[1589]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1397]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1398]_i_1 
       (.I0(\out[1526]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[417] ),
        .I2(\f_permutation_l_/out_reg_n_0_[40] ),
        .I3(\out[1462]_i_3_n_0 ),
        .I4(\out[1590]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1398]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1399]_i_1 
       (.I0(\out[1527]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[418] ),
        .I2(\f_permutation_l_/out_reg_n_0_[41] ),
        .I3(\out[1463]_i_3_n_0 ),
        .I4(\out[1591]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1399]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[139]_i_1 
       (.I0(\out[1458]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[676] ),
        .I2(\out[139]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[201] ),
        .I4(\out[1589]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [139]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[139]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[610] ),
        .I1(\f_permutation_l_/round_in [1505]),
        .I2(\out[1548]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[139]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[13]_i_1 
       (.I0(\out[1591]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[203] ),
        .I2(\out[269]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1046]),
        .I4(\out[1515]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1400]_i_1 
       (.I0(\out[1528]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[419] ),
        .I2(\f_permutation_l_/out_reg_n_0_[42] ),
        .I3(\out[1464]_i_3_n_0 ),
        .I4(\out[1592]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1400]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1401]_i_1 
       (.I0(\out[1529]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[420] ),
        .I2(\f_permutation_l_/out_reg_n_0_[43] ),
        .I3(\out[1465]_i_3_n_0 ),
        .I4(\out[1593]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1401]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1402]_i_1 
       (.I0(\out[1530]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[421] ),
        .I2(\f_permutation_l_/out_reg_n_0_[44] ),
        .I3(\out[1466]_i_3_n_0 ),
        .I4(\out[1594]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1402]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1403]_i_1 
       (.I0(\out[1531]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[422] ),
        .I2(\f_permutation_l_/out_reg_n_0_[45] ),
        .I3(\out[1467]_i_3_n_0 ),
        .I4(\out[1595]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1403]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1404]_i_1 
       (.I0(\out[1532]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[423] ),
        .I2(\f_permutation_l_/out_reg_n_0_[46] ),
        .I3(\out[1468]_i_3_n_0 ),
        .I4(\out[1596]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1404]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1405]_i_1 
       (.I0(\out[1533]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[424] ),
        .I2(\f_permutation_l_/out_reg_n_0_[47] ),
        .I3(\out[1469]_i_3_n_0 ),
        .I4(\out[1597]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1405]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1406]_i_1 
       (.I0(\out[1534]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[425] ),
        .I2(\f_permutation_l_/out_reg_n_0_[48] ),
        .I3(\out[1470]_i_3_n_0 ),
        .I4(\out[1598]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1406]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[1407]_i_1 
       (.I0(\out[1535]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[426] ),
        .I2(\f_permutation_l_/out_reg_n_0_[49] ),
        .I3(\out[1471]_i_3_n_0 ),
        .I4(\out[1599]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [1407]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1408]_i_1 
       (.I0(\out[1472]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[789] ),
        .I2(\out[1408]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[50] ),
        .I4(\out[1408]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1408]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1408]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[427] ),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[1408]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1408]_i_3 
       (.I0(\out[1566]_i_10_n_0 ),
        .I1(padder_out_1[330]),
        .I2(out[266]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1585]),
        .I5(\out[1565]_i_6_n_0 ),
        .O(\out[1408]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1409]_i_1 
       (.I0(\out[1537]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[790] ),
        .I2(\out[1409]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[51] ),
        .I4(\out[1409]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1409]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1409]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[428] ),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[1409]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1409]_i_3 
       (.I0(\out[1567]_i_11_n_0 ),
        .I1(padder_out_1[331]),
        .I2(out[267]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1586]),
        .I5(\out[1566]_i_6_n_0 ),
        .O(\out[1409]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[140]_i_1 
       (.I0(\out[1459]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[677] ),
        .I2(\out[140]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[202] ),
        .I4(\out[1590]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [140]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[140]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[611] ),
        .I1(\f_permutation_l_/round_in [1506]),
        .I2(\out[1549]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[140]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1410]_i_1 
       (.I0(\out[1538]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[791] ),
        .I2(\out[1410]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[52] ),
        .I4(\out[1410]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1410]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1410]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[429] ),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[1410]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1410]_i_3 
       (.I0(\out[1568]_i_10_n_0 ),
        .I1(padder_out_1[332]),
        .I2(out[268]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1587]),
        .I5(\out[1567]_i_9_n_0 ),
        .O(\out[1410]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[1411]_i_1 
       (.I0(\out[1539]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[430] ),
        .I2(\out[1475]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[53] ),
        .I4(\out[1411]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1411]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1411]_i_2 
       (.I0(\out[1569]_i_10_n_0 ),
        .I1(padder_out_1[333]),
        .I2(out[269]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1588]),
        .I5(\out[1568]_i_6_n_0 ),
        .O(\out[1411]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1412]_i_1 
       (.I0(\out[1540]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[793] ),
        .I2(\out[1412]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[54] ),
        .I4(\out[1412]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1412]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1412]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[431] ),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[1412]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1412]_i_3 
       (.I0(\out[1570]_i_10_n_0 ),
        .I1(padder_out_1[334]),
        .I2(out[270]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1589]),
        .I5(\out[1569]_i_6_n_0 ),
        .O(\out[1412]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1413]_i_1 
       (.I0(\out[1541]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[794] ),
        .I2(\out[1413]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[55] ),
        .I4(\out[1413]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1413]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1413]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[432] ),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[1413]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1413]_i_3 
       (.I0(\out[1571]_i_10_n_0 ),
        .I1(padder_out_1[335]),
        .I2(out[271]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1590]),
        .I5(\out[1570]_i_6_n_0 ),
        .O(\out[1413]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1414]_i_1 
       (.I0(\out[1542]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[795] ),
        .I2(\out[1414]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[56] ),
        .I4(\out[1414]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1414]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1414]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[433] ),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[1414]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1414]_i_3 
       (.I0(\out[1572]_i_10_n_0 ),
        .I1(padder_out_1[320]),
        .I2(out[256]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1591]),
        .I5(\out[1571]_i_6_n_0 ),
        .O(\out[1414]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1415]_i_1 
       (.I0(\out[1543]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[796] ),
        .I2(\out[1415]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[57] ),
        .I4(\out[1415]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1415]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1415]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[434] ),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[1415]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1415]_i_3 
       (.I0(\out[1573]_i_10_n_0 ),
        .I1(padder_out_1[321]),
        .I2(out[257]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1592]),
        .I5(\out[1572]_i_6_n_0 ),
        .O(\out[1415]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1415]_i_4 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1415]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1416]_i_1 
       (.I0(\out[1544]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[797] ),
        .I2(\out[1416]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[58] ),
        .I4(\out[1416]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1416]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1416]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[435] ),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[1416]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1416]_i_3 
       (.I0(\out[1574]_i_10_n_0 ),
        .I1(padder_out_1[322]),
        .I2(out[258]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1593]),
        .I5(\out[1573]_i_6_n_0 ),
        .O(\out[1416]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1417]_i_1 
       (.I0(\out[1545]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[798] ),
        .I2(\out[1417]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[59] ),
        .I4(\out[1417]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1417]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1417]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[436] ),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[1417]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1417]_i_3 
       (.I0(\out[1575]_i_10_n_0 ),
        .I1(padder_out_1[323]),
        .I2(out[259]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1594]),
        .I5(\out[1574]_i_6_n_0 ),
        .O(\out[1417]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1418]_i_1 
       (.I0(\out[1546]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[799] ),
        .I2(\out[1418]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[60] ),
        .I4(\out[1418]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1418]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1418]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[437] ),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[1418]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1418]_i_3 
       (.I0(\out[1576]_i_10_n_0 ),
        .I1(padder_out_1[324]),
        .I2(out[260]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1595]),
        .I5(\out[1575]_i_6_n_0 ),
        .O(\out[1418]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1419]_i_1 
       (.I0(\out[1547]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[800] ),
        .I2(\out[1419]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[61] ),
        .I4(\out[1419]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1419]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1419]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[438] ),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[1419]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1419]_i_3 
       (.I0(\out[1577]_i_10_n_0 ),
        .I1(padder_out_1[325]),
        .I2(out[261]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1596]),
        .I5(\out[1576]_i_6_n_0 ),
        .O(\out[1419]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[141]_i_1 
       (.I0(\out[1460]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[678] ),
        .I2(\out[141]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[203] ),
        .I4(\out[1591]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [141]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[141]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[612] ),
        .I1(\f_permutation_l_/round_in [1507]),
        .I2(\out[1550]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[141]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1420]_i_1 
       (.I0(\out[1548]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[801] ),
        .I2(\out[1420]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[62] ),
        .I4(\out[1420]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1420]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1420]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[439] ),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[1420]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1420]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[262]),
        .I2(padder_out_1[326]),
        .I3(\out[1578]_i_9_n_0 ),
        .I4(\out[1577]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1597]),
        .O(\out[1420]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1421]_i_1 
       (.I0(\out[1549]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[802] ),
        .I2(\out[1421]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[63] ),
        .I4(\out[1421]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1421]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1421]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[440] ),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[1421]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1421]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[263]),
        .I2(padder_out_1[327]),
        .I3(\out[1579]_i_10_n_0 ),
        .I4(\out[1578]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1598]),
        .O(\out[1421]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1422]_i_1 
       (.I0(\out[1550]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[803] ),
        .I2(\out[1422]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_ ),
        .I4(\out[1422]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1422]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1422]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[441] ),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[1422]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1422]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[312]),
        .I2(padder_out_1[376]),
        .I3(\out[1580]_i_9_n_0 ),
        .I4(\out[1579]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1599]),
        .O(\out[1422]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1423]_i_1 
       (.I0(\out[1551]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[804] ),
        .I2(\out[1423]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1] ),
        .I4(\out[1423]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1423]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1423]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[442] ),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[1423]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1423]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[313]),
        .I2(padder_out_1[377]),
        .I3(\out[1581]_i_9_n_0 ),
        .I4(\out[1580]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1536]),
        .O(\out[1423]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1424]_i_1 
       (.I0(\out[1552]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[805] ),
        .I2(\out[1424]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[2] ),
        .I4(\out[1424]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1424]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1424]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[443] ),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[1424]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1424]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[314]),
        .I2(padder_out_1[378]),
        .I3(\out[1582]_i_9_n_0 ),
        .I4(\out[1581]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1537]),
        .O(\out[1424]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1425]_i_1 
       (.I0(\out[1553]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[806] ),
        .I2(\out[1425]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[3] ),
        .I4(\out[1425]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1425]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1425]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[444] ),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[1425]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1425]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[315]),
        .I2(padder_out_1[379]),
        .I3(\out[1583]_i_9_n_0 ),
        .I4(\out[1582]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1538]),
        .O(\out[1425]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1426]_i_1 
       (.I0(\out[1554]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[807] ),
        .I2(\out[1426]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[4] ),
        .I4(\out[1426]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1426]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1426]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[445] ),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[1426]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1426]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[316]),
        .I2(padder_out_1[380]),
        .I3(\out[1584]_i_9_n_0 ),
        .I4(\out[1583]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1539]),
        .O(\out[1426]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1427]_i_1 
       (.I0(\out[1555]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[808] ),
        .I2(\out[1427]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[5] ),
        .I4(\out[1427]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1427]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1427]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[446] ),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[1427]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1427]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[317]),
        .I2(padder_out_1[381]),
        .I3(\out[1585]_i_9_n_0 ),
        .I4(\out[1584]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1540]),
        .O(\out[1427]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1428]_i_1 
       (.I0(\out[1556]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[809] ),
        .I2(\out[1428]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[6] ),
        .I4(\out[1428]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1428]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1428]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[447] ),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[1428]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1428]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[318]),
        .I2(padder_out_1[382]),
        .I3(\out[1586]_i_9_n_0 ),
        .I4(\out[1585]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1541]),
        .O(\out[1428]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1429]_i_1 
       (.I0(\out[1557]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[810] ),
        .I2(\out[1429]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[7] ),
        .I4(\out[1429]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1429]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1429]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[384] ),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[1429]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1429]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[319]),
        .I2(padder_out_1[383]),
        .I3(\out[1587]_i_9_n_0 ),
        .I4(\out[1586]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1542]),
        .O(\out[1429]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[142]_i_1 
       (.I0(\out[1461]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[679] ),
        .I2(\out[142]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[204] ),
        .I4(\out[1592]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [142]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[142]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[613] ),
        .I1(\f_permutation_l_/round_in [1508]),
        .I2(\out[1551]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[142]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1430]_i_1 
       (.I0(\out[1558]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[811] ),
        .I2(\out[1430]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[8] ),
        .I4(\out[1430]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1430]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1430]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[385] ),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1409]),
        .I4(\out[1582]_i_7_n_0 ),
        .O(\out[1430]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1430]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[304]),
        .I2(padder_out_1[368]),
        .I3(\out[1588]_i_9_n_0 ),
        .I4(\out[1587]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1543]),
        .O(\out[1430]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1431]_i_1 
       (.I0(\out[1559]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[812] ),
        .I2(\out[1431]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[9] ),
        .I4(\out[1431]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1431]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1431]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[386] ),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1410]),
        .I4(\out[1583]_i_7_n_0 ),
        .O(\out[1431]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1431]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[305]),
        .I2(padder_out_1[369]),
        .I3(\out[1589]_i_9_n_0 ),
        .I4(\out[1588]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1544]),
        .O(\out[1431]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1432]_i_1 
       (.I0(\out[1560]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[813] ),
        .I2(\out[1432]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[10] ),
        .I4(\out[1432]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1432]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1432]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[387] ),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1411]),
        .I4(\out[1584]_i_7_n_0 ),
        .O(\out[1432]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1432]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[306]),
        .I2(padder_out_1[370]),
        .I3(\out[1590]_i_9_n_0 ),
        .I4(\out[1589]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1545]),
        .O(\out[1432]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1433]_i_1 
       (.I0(\out[1561]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[814] ),
        .I2(\out[1433]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[11] ),
        .I4(\out[1433]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1433]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1433]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[388] ),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1412]),
        .I4(\out[1585]_i_7_n_0 ),
        .O(\out[1433]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1433]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[307]),
        .I2(padder_out_1[371]),
        .I3(\out[1591]_i_9_n_0 ),
        .I4(\out[1590]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1546]),
        .O(\out[1433]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1434]_i_1 
       (.I0(\out[1562]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[815] ),
        .I2(\out[1434]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[12] ),
        .I4(\out[1434]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1434]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1434]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[389] ),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1413]),
        .I4(\out[1586]_i_7_n_0 ),
        .O(\out[1434]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1434]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[308]),
        .I2(padder_out_1[372]),
        .I3(\out[1592]_i_9_n_0 ),
        .I4(\out[1591]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1547]),
        .O(\out[1434]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1435]_i_1 
       (.I0(\out[1563]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[816] ),
        .I2(\out[1435]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[13] ),
        .I4(\out[1435]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1435]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1435]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[390] ),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1414]),
        .I4(\out[1587]_i_7_n_0 ),
        .O(\out[1435]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1435]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[309]),
        .I2(padder_out_1[373]),
        .I3(\out[1593]_i_9_n_0 ),
        .I4(\out[1592]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1548]),
        .O(\out[1435]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1436]_i_1 
       (.I0(\out[1564]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[817] ),
        .I2(\out[1436]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[14] ),
        .I4(\out[1436]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1436]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1436]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[391] ),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1415]),
        .I4(\out[1588]_i_7_n_0 ),
        .O(\out[1436]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1436]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[310]),
        .I2(padder_out_1[374]),
        .I3(\out[1594]_i_9_n_0 ),
        .I4(\out[1593]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1549]),
        .O(\out[1436]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1437]_i_1 
       (.I0(\out[1565]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[818] ),
        .I2(\out[1437]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[15] ),
        .I4(\out[1437]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1437]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1437]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[392] ),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1416]),
        .I4(\out[1589]_i_7_n_0 ),
        .O(\out[1437]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1437]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[311]),
        .I2(padder_out_1[375]),
        .I3(\out[1595]_i_9_n_0 ),
        .I4(\out[1594]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1550]),
        .O(\out[1437]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1438]_i_1 
       (.I0(\out[1566]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[819] ),
        .I2(\out[1438]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[16] ),
        .I4(\out[1438]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1438]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1438]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[393] ),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1417]),
        .I4(\out[1590]_i_7_n_0 ),
        .O(\out[1438]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1438]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[296]),
        .I2(padder_out_1[360]),
        .I3(\out[1596]_i_9_n_0 ),
        .I4(\out[1595]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1551]),
        .O(\out[1438]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1439]_i_1 
       (.I0(\out[1567]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[820] ),
        .I2(\out[1439]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[17] ),
        .I4(\out[1439]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1439]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1439]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[394] ),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1418]),
        .I4(\out[1591]_i_7_n_0 ),
        .O(\out[1439]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1439]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[297]),
        .I2(padder_out_1[361]),
        .I3(\out[1597]_i_9_n_0 ),
        .I4(\out[1596]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1552]),
        .O(\out[1439]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[143]_i_1 
       (.I0(\out[1462]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[680] ),
        .I2(\out[143]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[205] ),
        .I4(\out[1593]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [143]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[143]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[614] ),
        .I1(\f_permutation_l_/round_in [1509]),
        .I2(\out[1552]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[143]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1440]_i_1 
       (.I0(\out[1568]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[821] ),
        .I2(\out[1440]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[18] ),
        .I4(\out[1440]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1440]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1440]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[395] ),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1419]),
        .I4(\out[1592]_i_7_n_0 ),
        .O(\out[1440]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1440]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[298]),
        .I2(padder_out_1[362]),
        .I3(\out[1598]_i_9_n_0 ),
        .I4(\out[1597]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1553]),
        .O(\out[1440]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1441]_i_1 
       (.I0(\out[1569]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[822] ),
        .I2(\out[1441]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[19] ),
        .I4(\out[1441]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1441]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1441]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[396] ),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1420]),
        .I4(\out[1593]_i_7_n_0 ),
        .O(\out[1441]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1441]_i_3 
       (.I0(\out[1415]_i_4_n_0 ),
        .I1(out[299]),
        .I2(padder_out_1[363]),
        .I3(\out[1599]_i_9_n_0 ),
        .I4(\out[1598]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1554]),
        .O(\out[1441]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[1442]_i_1 
       (.I0(\out[1570]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[823] ),
        .I2(\out[1442]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[20] ),
        .I4(\out[1442]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1442]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1442]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[397] ),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1421]),
        .I4(\out[1594]_i_7_n_0 ),
        .O(\out[1442]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1442]_i_3 
       (.I0(\out[1599]_i_8_n_0 ),
        .I1(padder_out_1[555]),
        .I2(out[491]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1536]_i_12_n_0 ),
        .I5(\f_permutation_l_/round_in [1364]),
        .O(\out[1442]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1443]_i_1 
       (.I0(\out[1571]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[824] ),
        .I2(\out[1443]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[21] ),
        .I4(\out[1443]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1443]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1443]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[398] ),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1422]),
        .I4(\out[1595]_i_7_n_0 ),
        .O(\out[1443]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1443]_i_3 
       (.I0(\out[1537]_i_11_n_0 ),
        .I1(padder_out_1[365]),
        .I2(out[301]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1556]),
        .I5(\out[1536]_i_10_n_0 ),
        .O(\out[1443]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1444]_i_1 
       (.I0(\out[1572]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[825] ),
        .I2(\out[1444]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[22] ),
        .I4(\out[1444]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1444]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1444]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[399] ),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1423]),
        .I4(\out[1596]_i_7_n_0 ),
        .O(\out[1444]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1444]_i_3 
       (.I0(\out[1538]_i_10_n_0 ),
        .I1(padder_out_1[366]),
        .I2(out[302]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1557]),
        .I5(\out[1537]_i_9_n_0 ),
        .O(\out[1444]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1445]_i_1 
       (.I0(\out[1573]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[826] ),
        .I2(\out[1445]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[23] ),
        .I4(\out[1445]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1445]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1445]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[400] ),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1424]),
        .I4(\out[1597]_i_7_n_0 ),
        .O(\out[1445]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1445]_i_3 
       (.I0(\out[1447]_i_4_n_0 ),
        .I1(out[303]),
        .I2(padder_out_1[367]),
        .I3(\out[1539]_i_12_n_0 ),
        .I4(\out[1538]_i_6_n_0 ),
        .I5(\f_permutation_l_/round_in [1558]),
        .O(\out[1445]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1446]_i_1 
       (.I0(\out[1574]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[827] ),
        .I2(\out[1446]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[24] ),
        .I4(\out[1446]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1446]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1446]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[401] ),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1425]),
        .I4(\out[1598]_i_7_n_0 ),
        .O(\out[1446]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1446]_i_3 
       (.I0(\out[1540]_i_10_n_0 ),
        .I1(padder_out_1[352]),
        .I2(out[288]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1559]),
        .I5(\out[1539]_i_8_n_0 ),
        .O(\out[1446]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1447]_i_1 
       (.I0(\out[1575]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[828] ),
        .I2(\out[1447]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[25] ),
        .I4(\out[1447]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1447]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1447]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[402] ),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\out[1599]_i_7_n_0 ),
        .I4(\f_permutation_l_/round_in [1426]),
        .O(\out[1447]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1447]_i_3 
       (.I0(\out[1541]_i_10_n_0 ),
        .I1(padder_out_1[353]),
        .I2(out[289]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1560]),
        .I5(\out[1540]_i_6_n_0 ),
        .O(\out[1447]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1447]_i_4 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1447]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1448]_i_1 
       (.I0(\out[1576]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[829] ),
        .I2(\out[1448]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[26] ),
        .I4(\out[1448]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1448]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1448]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[403] ),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\out[1554]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1298]),
        .O(\out[1448]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1448]_i_3 
       (.I0(\out[1542]_i_12_n_0 ),
        .I1(padder_out_1[354]),
        .I2(out[290]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1561]),
        .I5(\out[1541]_i_6_n_0 ),
        .O(\out[1448]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[1449]_i_1 
       (.I0(\out[1577]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[830] ),
        .I2(\out[1449]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[27] ),
        .I4(\out[1449]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1449]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1449]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[404] ),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\out[1555]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1299]),
        .O(\out[1449]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1449]_i_3 
       (.I0(\out[1543]_i_13_n_0 ),
        .I1(padder_out_1[355]),
        .I2(out[291]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1562]),
        .I5(\out[1542]_i_7_n_0 ),
        .O(\out[1449]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[144]_i_1 
       (.I0(\out[1463]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[681] ),
        .I2(\out[144]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[206] ),
        .I4(\out[1594]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [144]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[144]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[615] ),
        .I1(\f_permutation_l_/round_in [1510]),
        .I2(\out[1553]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[144]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1450]_i_1 
       (.I0(\out[1578]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[831] ),
        .I2(\out[1450]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[28] ),
        .I4(\out[1450]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1450]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1450]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[405] ),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\out[1556]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1300]),
        .O(\out[1450]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1450]_i_3 
       (.I0(\out[1544]_i_10_n_0 ),
        .I1(padder_out_1[356]),
        .I2(out[292]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1563]),
        .I5(\out[1543]_i_10_n_0 ),
        .O(\out[1450]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1451]_i_1 
       (.I0(\out[1579]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[768] ),
        .I2(\out[1451]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[29] ),
        .I4(\out[1451]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1451]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1451]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[406] ),
        .I1(\f_permutation_l_/round_in [1430]),
        .I2(\out[1539]_i_9_n_0 ),
        .I3(\out[1557]_i_13_n_0 ),
        .I4(\f_permutation_l_/round_in [1301]),
        .O(\out[1451]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1451]_i_3 
       (.I0(\out[1545]_i_10_n_0 ),
        .I1(padder_out_1[357]),
        .I2(out[293]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1564]),
        .I5(\out[1544]_i_6_n_0 ),
        .O(\out[1451]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1452]_i_1 
       (.I0(\out[1580]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[769] ),
        .I2(\out[1452]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[30] ),
        .I4(\out[1452]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1452]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1452]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[407] ),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[1452]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1452]_i_3 
       (.I0(\out[1546]_i_10_n_0 ),
        .I1(padder_out_1[358]),
        .I2(out[294]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1565]),
        .I5(\out[1545]_i_6_n_0 ),
        .O(\out[1452]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1453]_i_1 
       (.I0(\out[1581]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[770] ),
        .I2(\out[1453]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[31] ),
        .I4(\out[1453]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1453]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1453]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[408] ),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[1453]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1453]_i_3 
       (.I0(\out[1547]_i_10_n_0 ),
        .I1(padder_out_1[359]),
        .I2(out[295]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1566]),
        .I5(\out[1546]_i_6_n_0 ),
        .O(\out[1453]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1454]_i_1 
       (.I0(\out[1582]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[771] ),
        .I2(\out[1454]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[32] ),
        .I4(\out[1454]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1454]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1454]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[409] ),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[1454]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1454]_i_3 
       (.I0(\out[1548]_i_10_n_0 ),
        .I1(padder_out_1[344]),
        .I2(out[280]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1567]),
        .I5(\out[1547]_i_6_n_0 ),
        .O(\out[1454]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1455]_i_1 
       (.I0(\out[1583]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[772] ),
        .I2(\out[1455]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[33] ),
        .I4(\out[1455]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1455]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1455]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[410] ),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[1455]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1455]_i_3 
       (.I0(\out[1549]_i_10_n_0 ),
        .I1(padder_out_1[345]),
        .I2(out[281]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1568]),
        .I5(\out[1548]_i_6_n_0 ),
        .O(\out[1455]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1456]_i_1 
       (.I0(\out[1584]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[773] ),
        .I2(\out[1456]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[34] ),
        .I4(\out[1456]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1456]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1456]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[411] ),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[1456]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1456]_i_3 
       (.I0(\out[1550]_i_10_n_0 ),
        .I1(padder_out_1[346]),
        .I2(out[282]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1569]),
        .I5(\out[1549]_i_6_n_0 ),
        .O(\out[1456]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1457]_i_1 
       (.I0(\out[1585]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[774] ),
        .I2(\out[1457]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[35] ),
        .I4(\out[1457]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1457]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1457]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[412] ),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[1457]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1457]_i_3 
       (.I0(\out[1551]_i_11_n_0 ),
        .I1(padder_out_1[347]),
        .I2(out[283]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1570]),
        .I5(\out[1550]_i_6_n_0 ),
        .O(\out[1457]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1458]_i_1 
       (.I0(\out[1586]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[775] ),
        .I2(\out[1458]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[36] ),
        .I4(\out[1458]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1458]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1458]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[413] ),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[1458]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1458]_i_3 
       (.I0(\out[1552]_i_10_n_0 ),
        .I1(padder_out_1[348]),
        .I2(out[284]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1571]),
        .I5(\out[1551]_i_9_n_0 ),
        .O(\out[1458]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1459]_i_1 
       (.I0(\out[1587]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[776] ),
        .I2(\out[1459]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[37] ),
        .I4(\out[1459]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1459]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1459]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[414] ),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[1459]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1459]_i_3 
       (.I0(\out[1553]_i_10_n_0 ),
        .I1(padder_out_1[349]),
        .I2(out[285]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1572]),
        .I5(\out[1552]_i_6_n_0 ),
        .O(\out[1459]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[145]_i_1 
       (.I0(\out[1464]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[682] ),
        .I2(\out[145]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[207] ),
        .I4(\out[1595]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [145]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[145]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[616] ),
        .I1(\f_permutation_l_/round_in [1511]),
        .I2(\out[1554]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[145]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1460]_i_1 
       (.I0(\out[1588]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[777] ),
        .I2(\out[1460]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[38] ),
        .I4(\out[1460]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1460]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1460]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[415] ),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[1460]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1460]_i_3 
       (.I0(\out[1554]_i_10_n_0 ),
        .I1(padder_out_1[350]),
        .I2(out[286]),
        .I3(\out[1447]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1573]),
        .I5(\out[1553]_i_6_n_0 ),
        .O(\out[1460]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1461]_i_1 
       (.I0(\out[1589]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[778] ),
        .I2(\out[1461]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[39] ),
        .I4(\out[1461]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1461]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1461]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[416] ),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[1461]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1461]_i_3 
       (.I0(\out[1555]_i_10_n_0 ),
        .I1(padder_out_1[351]),
        .I2(out[287]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1574]),
        .I5(\out[1554]_i_6_n_0 ),
        .O(\out[1461]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1462]_i_1 
       (.I0(\out[1590]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[779] ),
        .I2(\out[1462]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[40] ),
        .I4(\out[1462]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1462]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1462]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[417] ),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[1462]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1462]_i_3 
       (.I0(\out[1556]_i_11_n_0 ),
        .I1(padder_out_1[336]),
        .I2(out[272]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1575]),
        .I5(\out[1555]_i_6_n_0 ),
        .O(\out[1462]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1463]_i_1 
       (.I0(\out[1591]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[780] ),
        .I2(\out[1463]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[41] ),
        .I4(\out[1463]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1463]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1463]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[418] ),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[1463]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1463]_i_3 
       (.I0(\out[1557]_i_10_n_0 ),
        .I1(padder_out_1[337]),
        .I2(out[273]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1576]),
        .I5(\out[1556]_i_6_n_0 ),
        .O(\out[1463]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1464]_i_1 
       (.I0(\out[1592]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[781] ),
        .I2(\out[1464]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[42] ),
        .I4(\out[1464]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1464]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1464]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[419] ),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[1464]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1464]_i_3 
       (.I0(\out[1558]_i_10_n_0 ),
        .I1(padder_out_1[338]),
        .I2(out[274]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1577]),
        .I5(\out[1557]_i_6_n_0 ),
        .O(\out[1464]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1465]_i_1 
       (.I0(\out[1593]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[782] ),
        .I2(\out[1465]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[43] ),
        .I4(\out[1465]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1465]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1465]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[420] ),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[1465]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1465]_i_3 
       (.I0(\out[1559]_i_10_n_0 ),
        .I1(padder_out_1[339]),
        .I2(out[275]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1578]),
        .I5(\out[1558]_i_6_n_0 ),
        .O(\out[1465]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1466]_i_1 
       (.I0(\out[1594]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[783] ),
        .I2(\out[1466]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[44] ),
        .I4(\out[1466]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1466]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1466]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[421] ),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[1466]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1466]_i_3 
       (.I0(\out[1560]_i_10_n_0 ),
        .I1(padder_out_1[340]),
        .I2(out[276]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1579]),
        .I5(\out[1559]_i_6_n_0 ),
        .O(\out[1466]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1467]_i_1 
       (.I0(\out[1595]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[784] ),
        .I2(\out[1467]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[45] ),
        .I4(\out[1467]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1467]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1467]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[422] ),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[1467]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1467]_i_3 
       (.I0(\out[1561]_i_10_n_0 ),
        .I1(padder_out_1[341]),
        .I2(out[277]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1580]),
        .I5(\out[1560]_i_6_n_0 ),
        .O(\out[1467]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1468]_i_1 
       (.I0(\out[1596]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[785] ),
        .I2(\out[1468]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[46] ),
        .I4(\out[1468]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1468]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1468]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[423] ),
        .I1(\f_permutation_l_/round_in [1447]),
        .I2(\out[1556]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[1468]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1468]_i_3 
       (.I0(\out[1562]_i_10_n_0 ),
        .I1(padder_out_1[342]),
        .I2(out[278]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1581]),
        .I5(\out[1561]_i_6_n_0 ),
        .O(\out[1468]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1469]_i_1 
       (.I0(\out[1597]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[786] ),
        .I2(\out[1469]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[47] ),
        .I4(\out[1469]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1469]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1469]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[424] ),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[1469]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1469]_i_3 
       (.I0(\out[1563]_i_10_n_0 ),
        .I1(padder_out_1[343]),
        .I2(out[279]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1582]),
        .I5(\out[1562]_i_6_n_0 ),
        .O(\out[1469]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[146]_i_1 
       (.I0(\out[1465]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[683] ),
        .I2(\out[146]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[208] ),
        .I4(\out[1596]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [146]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[146]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[617] ),
        .I1(\f_permutation_l_/round_in [1512]),
        .I2(\out[1555]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[146]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1470]_i_1 
       (.I0(\out[1598]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[787] ),
        .I2(\out[1470]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[48] ),
        .I4(\out[1470]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1470]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1470]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[425] ),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[1470]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1470]_i_3 
       (.I0(\out[1564]_i_10_n_0 ),
        .I1(padder_out_1[328]),
        .I2(out[264]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1583]),
        .I5(\out[1563]_i_6_n_0 ),
        .O(\out[1470]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[1471]_i_1 
       (.I0(\out[1599]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[788] ),
        .I2(\out[1471]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[49] ),
        .I4(\out[1471]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1471]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1471]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[426] ),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[1471]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1471]_i_3 
       (.I0(\out[1565]_i_10_n_0 ),
        .I1(padder_out_1[329]),
        .I2(out[265]),
        .I3(\out[1415]_i_4_n_0 ),
        .I4(\f_permutation_l_/round_in [1584]),
        .I5(\out[1564]_i_6_n_0 ),
        .O(\out[1471]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1472]_i_1 
       (.I0(\out[1536]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[789] ),
        .I2(\out[1472]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[427] ),
        .I4(\out[1472]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1472]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1472]_i_2 
       (.I0(\out[1536]_i_14_n_0 ),
        .I1(padder_out_1[493]),
        .I2(out[429]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1536]_i_12_n_0 ),
        .I5(\f_permutation_l_/round_in [1364]),
        .O(\out[1472]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1472]_i_3 
       (.I0(\out[1578]_i_14_n_0 ),
        .I1(padder_out_1[274]),
        .I2(out[210]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1560]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1451]),
        .O(\out[1472]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1473]_i_1 
       (.I0(\out[1537]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[790] ),
        .I2(\out[1537]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[428] ),
        .I4(\out[1473]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1473]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1473]_i_2 
       (.I0(\out[1579]_i_15_n_0 ),
        .I1(padder_out_1[275]),
        .I2(out[211]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1561]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1452]),
        .O(\out[1473]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1474]_i_1 
       (.I0(\out[1474]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[791] ),
        .I2(\out[1538]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[429] ),
        .I4(\out[1474]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1474]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1474]_i_2 
       (.I0(\f_permutation_l_/round_in [1174]),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1558]),
        .I4(\out[1538]_i_6_n_0 ),
        .O(\out[1474]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1474]_i_3 
       (.I0(\out[1580]_i_14_n_0 ),
        .I1(padder_out_1[276]),
        .I2(out[212]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1562]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1453]),
        .O(\out[1474]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1475]_i_1 
       (.I0(\out[1539]_i_3_n_0 ),
        .I1(\f_permutation_l_/round_in [1175]),
        .I2(\out[1539]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[430] ),
        .I4(\out[1475]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1475]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1475]_i_2 
       (.I0(\out[1581]_i_14_n_0 ),
        .I1(padder_out_1[277]),
        .I2(out[213]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1563]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1454]),
        .O(\out[1475]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1476]_i_1 
       (.I0(\out[1476]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[793] ),
        .I2(\out[1540]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[431] ),
        .I4(\out[1476]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1476]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1476]_i_2 
       (.I0(\f_permutation_l_/round_in [1176]),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1560]),
        .I4(\out[1540]_i_6_n_0 ),
        .O(\out[1476]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1476]_i_3 
       (.I0(\out[1582]_i_14_n_0 ),
        .I1(padder_out_1[278]),
        .I2(out[214]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1564]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1455]),
        .O(\out[1476]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1477]_i_1 
       (.I0(\out[1477]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[794] ),
        .I2(\out[1541]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[432] ),
        .I4(\out[1477]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1477]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1477]_i_2 
       (.I0(\f_permutation_l_/round_in [1177]),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1561]),
        .I4(\out[1541]_i_6_n_0 ),
        .O(\out[1477]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1477]_i_3 
       (.I0(\out[1583]_i_14_n_0 ),
        .I1(padder_out_1[279]),
        .I2(out[215]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1565]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1456]),
        .O(\out[1477]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1478]_i_1 
       (.I0(\out[1478]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[795] ),
        .I2(\out[1542]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[433] ),
        .I4(\out[1478]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1478]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1478]_i_2 
       (.I0(\f_permutation_l_/round_in [1178]),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1562]),
        .I4(\out[1542]_i_7_n_0 ),
        .O(\out[1478]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1478]_i_3 
       (.I0(\out[1584]_i_14_n_0 ),
        .I1(padder_out_1[264]),
        .I2(out[200]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1566]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1457]),
        .O(\out[1478]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1479]_i_1 
       (.I0(\out[1543]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[796] ),
        .I2(\out[1543]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[434] ),
        .I4(\out[1479]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1479]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1479]_i_2 
       (.I0(\out[1585]_i_14_n_0 ),
        .I1(padder_out_1[265]),
        .I2(out[201]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1567]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1458]),
        .O(\out[1479]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[147]_i_1 
       (.I0(\out[1466]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[684] ),
        .I2(\out[147]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[209] ),
        .I4(\out[1597]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [147]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[147]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[618] ),
        .I1(\f_permutation_l_/round_in [1513]),
        .I2(\out[1556]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[147]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1480]_i_1 
       (.I0(\out[1480]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[797] ),
        .I2(\out[1544]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[435] ),
        .I4(\out[1480]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1480]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1480]_i_2 
       (.I0(\f_permutation_l_/round_in [1180]),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1564]),
        .I4(\out[1544]_i_6_n_0 ),
        .O(\out[1480]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1480]_i_3 
       (.I0(\out[1586]_i_14_n_0 ),
        .I1(padder_out_1[266]),
        .I2(out[202]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1568]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1459]),
        .O(\out[1480]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1481]_i_1 
       (.I0(\out[1481]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[798] ),
        .I2(\out[1545]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[436] ),
        .I4(\out[1481]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1481]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1481]_i_2 
       (.I0(\f_permutation_l_/round_in [1181]),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1565]),
        .I4(\out[1545]_i_6_n_0 ),
        .O(\out[1481]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1481]_i_3 
       (.I0(\out[1587]_i_13_n_0 ),
        .I1(padder_out_1[267]),
        .I2(out[203]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1569]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1460]),
        .O(\out[1481]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1482]_i_1 
       (.I0(\out[1482]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[799] ),
        .I2(\out[1546]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[437] ),
        .I4(\out[1482]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1482]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1482]_i_2 
       (.I0(\f_permutation_l_/round_in [1182]),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1566]),
        .I4(\out[1546]_i_6_n_0 ),
        .O(\out[1482]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1482]_i_3 
       (.I0(\out[1588]_i_14_n_0 ),
        .I1(padder_out_1[268]),
        .I2(out[204]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1570]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1461]),
        .O(\out[1482]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1483]_i_1 
       (.I0(\out[1483]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[800] ),
        .I2(\out[1547]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[438] ),
        .I4(\out[1483]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1483]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1483]_i_2 
       (.I0(\f_permutation_l_/round_in [1183]),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1567]),
        .I4(\out[1547]_i_6_n_0 ),
        .O(\out[1483]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1483]_i_3 
       (.I0(\out[1589]_i_14_n_0 ),
        .I1(padder_out_1[269]),
        .I2(out[205]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1571]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1462]),
        .O(\out[1483]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1484]_i_1 
       (.I0(\out[1484]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[801] ),
        .I2(\out[1548]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[439] ),
        .I4(\out[1484]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1484]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1484]_i_2 
       (.I0(\f_permutation_l_/round_in [1184]),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1568]),
        .I4(\out[1548]_i_6_n_0 ),
        .O(\out[1484]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1484]_i_3 
       (.I0(\out[1590]_i_14_n_0 ),
        .I1(padder_out_1[270]),
        .I2(out[206]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1572]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1463]),
        .O(\out[1484]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1485]_i_1 
       (.I0(\out[1485]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[802] ),
        .I2(\out[1549]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[440] ),
        .I4(\out[1485]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1485]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1485]_i_2 
       (.I0(\f_permutation_l_/round_in [1185]),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1569]),
        .I4(\out[1549]_i_6_n_0 ),
        .O(\out[1485]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1485]_i_3 
       (.I0(\out[1591]_i_14_n_0 ),
        .I1(padder_out_1[271]),
        .I2(out[207]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1573]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1464]),
        .O(\out[1485]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1486]_i_1 
       (.I0(\out[1486]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[803] ),
        .I2(\out[1550]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[441] ),
        .I4(\out[1486]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1486]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1486]_i_2 
       (.I0(\f_permutation_l_/round_in [1186]),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1570]),
        .I4(\out[1550]_i_6_n_0 ),
        .O(\out[1486]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1486]_i_3 
       (.I0(\out[1592]_i_14_n_0 ),
        .I1(padder_out_1[256]),
        .I2(out[192]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1574]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1465]),
        .O(\out[1486]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1487]_i_1 
       (.I0(\out[1551]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[804] ),
        .I2(\out[1551]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[442] ),
        .I4(\out[1487]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1487]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1487]_i_2 
       (.I0(\out[1593]_i_14_n_0 ),
        .I1(padder_out_1[257]),
        .I2(out[193]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1575]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1466]),
        .O(\out[1487]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1488]_i_1 
       (.I0(\out[1488]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[805] ),
        .I2(\out[1552]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[443] ),
        .I4(\out[1488]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1488]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1488]_i_2 
       (.I0(\f_permutation_l_/round_in [1188]),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1572]),
        .I4(\out[1552]_i_6_n_0 ),
        .O(\out[1488]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1488]_i_3 
       (.I0(\out[1594]_i_14_n_0 ),
        .I1(padder_out_1[258]),
        .I2(out[194]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1576]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1467]),
        .O(\out[1488]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1489]_i_1 
       (.I0(\out[1489]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[806] ),
        .I2(\out[1553]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[444] ),
        .I4(\out[1489]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1489]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1489]_i_2 
       (.I0(\f_permutation_l_/round_in [1189]),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1573]),
        .I4(\out[1553]_i_6_n_0 ),
        .O(\out[1489]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1489]_i_3 
       (.I0(\out[1595]_i_14_n_0 ),
        .I1(padder_out_1[259]),
        .I2(out[195]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1577]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1468]),
        .O(\out[1489]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[148]_i_1 
       (.I0(\out[1467]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[685] ),
        .I2(\out[148]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[210] ),
        .I4(\out[1598]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [148]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[148]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[619] ),
        .I1(\f_permutation_l_/round_in [1514]),
        .I2(\out[1557]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[148]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1490]_i_1 
       (.I0(\out[1490]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[807] ),
        .I2(\out[1554]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[445] ),
        .I4(\out[1490]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1490]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1490]_i_2 
       (.I0(\f_permutation_l_/round_in [1190]),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1574]),
        .I4(\out[1554]_i_6_n_0 ),
        .O(\out[1490]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1490]_i_3 
       (.I0(\out[1596]_i_14_n_0 ),
        .I1(padder_out_1[260]),
        .I2(out[196]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1578]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1469]),
        .O(\out[1490]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1491]_i_1 
       (.I0(\out[1491]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[808] ),
        .I2(\out[1555]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[446] ),
        .I4(\out[1491]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1491]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1491]_i_2 
       (.I0(\f_permutation_l_/round_in [1191]),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1575]),
        .I4(\out[1555]_i_6_n_0 ),
        .O(\out[1491]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1491]_i_3 
       (.I0(\out[1597]_i_14_n_0 ),
        .I1(padder_out_1[261]),
        .I2(out[197]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1579]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1470]),
        .O(\out[1491]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1492]_i_1 
       (.I0(\out[1492]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[809] ),
        .I2(\out[1556]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[447] ),
        .I4(\out[1492]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1492]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1492]_i_2 
       (.I0(\f_permutation_l_/round_in [1192]),
        .I1(\f_permutation_l_/round_in [1447]),
        .I2(\out[1556]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1576]),
        .I4(\out[1556]_i_6_n_0 ),
        .O(\out[1492]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1492]_i_3 
       (.I0(\out[1598]_i_14_n_0 ),
        .I1(padder_out_1[262]),
        .I2(out[198]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1580]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1471]),
        .O(\out[1492]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1493]_i_1 
       (.I0(\out[1493]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[810] ),
        .I2(\out[1557]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[384] ),
        .I4(\out[1493]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1493]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1493]_i_2 
       (.I0(\f_permutation_l_/round_in [1193]),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1577]),
        .I4(\out[1557]_i_6_n_0 ),
        .O(\out[1493]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1493]_i_3 
       (.I0(\out[1599]_i_14_n_0 ),
        .I1(padder_out_1[263]),
        .I2(out[199]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1581]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1408]),
        .O(\out[1493]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1494]_i_1 
       (.I0(\out[1494]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[811] ),
        .I2(\out[1558]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[385] ),
        .I4(\out[1494]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1494]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1494]_i_2 
       (.I0(\f_permutation_l_/round_in [1194]),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1578]),
        .I4(\out[1558]_i_6_n_0 ),
        .O(\out[1494]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1494]_i_3 
       (.I0(\out[1582]_i_7_n_0 ),
        .I1(padder_out_1[441]),
        .I2(out[377]),
        .I3(\i[0]_i_1__0_n_0 ),
        .I4(\out[1536]_i_17_n_0 ),
        .I5(\f_permutation_l_/round_in [1280]),
        .O(\out[1494]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1495]_i_1 
       (.I0(\out[1495]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[812] ),
        .I2(\out[1559]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[386] ),
        .I4(\out[1495]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1495]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1495]_i_2 
       (.I0(\f_permutation_l_/round_in [1195]),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1579]),
        .I4(\out[1559]_i_6_n_0 ),
        .O(\out[1495]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1495]_i_3 
       (.I0(\out[1583]_i_7_n_0 ),
        .I1(padder_out_1[442]),
        .I2(out[378]),
        .I3(\i[0]_i_1__0_n_0 ),
        .I4(\out[1537]_i_15_n_0 ),
        .I5(\f_permutation_l_/round_in [1281]),
        .O(\out[1495]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1496]_i_1 
       (.I0(\out[1496]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[813] ),
        .I2(\out[1560]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[387] ),
        .I4(\out[1496]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1496]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1496]_i_2 
       (.I0(\f_permutation_l_/round_in [1196]),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1580]),
        .I4(\out[1560]_i_6_n_0 ),
        .O(\out[1496]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1496]_i_3 
       (.I0(\out[1584]_i_7_n_0 ),
        .I1(padder_out_1[443]),
        .I2(out[379]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1538]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1282]),
        .O(\out[1496]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1497]_i_1 
       (.I0(\out[1497]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[814] ),
        .I2(\out[1561]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[388] ),
        .I4(\out[1497]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1497]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1497]_i_2 
       (.I0(\f_permutation_l_/round_in [1197]),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1581]),
        .I4(\out[1561]_i_6_n_0 ),
        .O(\out[1497]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1497]_i_3 
       (.I0(\out[1585]_i_7_n_0 ),
        .I1(padder_out_1[444]),
        .I2(out[380]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1539]_i_16_n_0 ),
        .I5(\f_permutation_l_/round_in [1283]),
        .O(\out[1497]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1498]_i_1 
       (.I0(\out[1498]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[815] ),
        .I2(\out[1562]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[389] ),
        .I4(\out[1498]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1498]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1498]_i_2 
       (.I0(\f_permutation_l_/round_in [1198]),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1582]),
        .I4(\out[1562]_i_6_n_0 ),
        .O(\out[1498]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1498]_i_3 
       (.I0(\out[1586]_i_7_n_0 ),
        .I1(padder_out_1[445]),
        .I2(out[381]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1540]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1284]),
        .O(\out[1498]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1499]_i_1 
       (.I0(\out[1499]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[816] ),
        .I2(\out[1563]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[390] ),
        .I4(\out[1499]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1499]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1499]_i_2 
       (.I0(\f_permutation_l_/round_in [1199]),
        .I1(\f_permutation_l_/round_in [1454]),
        .I2(\out[1563]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1583]),
        .I4(\out[1563]_i_6_n_0 ),
        .O(\out[1499]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1499]_i_3 
       (.I0(\out[1587]_i_7_n_0 ),
        .I1(padder_out_1[446]),
        .I2(out[382]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1541]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1285]),
        .O(\out[1499]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[149]_i_1 
       (.I0(\out[1468]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[686] ),
        .I2(\out[149]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[211] ),
        .I4(\out[1343]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [149]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[149]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[620] ),
        .I1(\f_permutation_l_/round_in [1515]),
        .I2(\out[1558]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[149]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[14]_i_1 
       (.I0(\out[1592]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[204] ),
        .I2(\out[270]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1047]),
        .I4(\out[1516]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1500]_i_1 
       (.I0(\out[1500]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[817] ),
        .I2(\out[1564]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[391] ),
        .I4(\out[1500]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1500]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1500]_i_2 
       (.I0(\f_permutation_l_/round_in [1200]),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1584]),
        .I4(\out[1564]_i_6_n_0 ),
        .O(\out[1500]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1500]_i_3 
       (.I0(\out[1588]_i_7_n_0 ),
        .I1(padder_out_1[447]),
        .I2(out[383]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1542]_i_16_n_0 ),
        .I5(\f_permutation_l_/round_in [1286]),
        .O(\out[1500]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1501]_i_1 
       (.I0(\out[1501]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[818] ),
        .I2(\out[1565]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[392] ),
        .I4(\out[1501]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1501]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1501]_i_2 
       (.I0(\f_permutation_l_/round_in [1201]),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1585]),
        .I4(\out[1565]_i_6_n_0 ),
        .O(\out[1501]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1501]_i_3 
       (.I0(\out[1589]_i_7_n_0 ),
        .I1(padder_out_1[432]),
        .I2(out[368]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1543]_i_17_n_0 ),
        .I5(\f_permutation_l_/round_in [1287]),
        .O(\out[1501]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1502]_i_1 
       (.I0(\out[1502]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[819] ),
        .I2(\out[1566]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[393] ),
        .I4(\out[1502]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1502]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1502]_i_2 
       (.I0(\f_permutation_l_/round_in [1202]),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1586]),
        .I4(\out[1566]_i_6_n_0 ),
        .O(\out[1502]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1502]_i_3 
       (.I0(\out[1590]_i_7_n_0 ),
        .I1(padder_out_1[433]),
        .I2(out[369]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1544]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1288]),
        .O(\out[1502]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1503]_i_1 
       (.I0(\out[1567]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[820] ),
        .I2(\out[1567]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[394] ),
        .I4(\out[1503]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1503]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1503]_i_2 
       (.I0(\out[1591]_i_7_n_0 ),
        .I1(padder_out_1[434]),
        .I2(out[370]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1545]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1289]),
        .O(\out[1503]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1504]_i_1 
       (.I0(\out[1504]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[821] ),
        .I2(\out[1568]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[395] ),
        .I4(\out[1504]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1504]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1504]_i_2 
       (.I0(\f_permutation_l_/round_in [1204]),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1588]),
        .I4(\out[1568]_i_6_n_0 ),
        .O(\out[1504]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1504]_i_3 
       (.I0(\out[1592]_i_7_n_0 ),
        .I1(padder_out_1[435]),
        .I2(out[371]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1546]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1290]),
        .O(\out[1504]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1505]_i_1 
       (.I0(\out[1505]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[822] ),
        .I2(\out[1569]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[396] ),
        .I4(\out[1505]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1505]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1505]_i_2 
       (.I0(\f_permutation_l_/round_in [1205]),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1589]),
        .I4(\out[1569]_i_6_n_0 ),
        .O(\out[1505]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1505]_i_3 
       (.I0(\out[1593]_i_7_n_0 ),
        .I1(padder_out_1[436]),
        .I2(out[372]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1547]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1291]),
        .O(\out[1505]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1506]_i_1 
       (.I0(\out[1506]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[823] ),
        .I2(\out[1570]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[397] ),
        .I4(\out[1506]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1506]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1506]_i_2 
       (.I0(\f_permutation_l_/round_in [1206]),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1590]),
        .I4(\out[1570]_i_6_n_0 ),
        .O(\out[1506]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1506]_i_3 
       (.I0(\out[1594]_i_7_n_0 ),
        .I1(padder_out_1[437]),
        .I2(out[373]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1548]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1292]),
        .O(\out[1506]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1507]_i_1 
       (.I0(\out[1507]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[824] ),
        .I2(\out[1571]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[398] ),
        .I4(\out[1507]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1507]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1507]_i_2 
       (.I0(\f_permutation_l_/round_in [1207]),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1591]),
        .I4(\out[1571]_i_6_n_0 ),
        .O(\out[1507]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1507]_i_3 
       (.I0(\out[1595]_i_7_n_0 ),
        .I1(padder_out_1[438]),
        .I2(out[374]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1549]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1293]),
        .O(\out[1507]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1508]_i_1 
       (.I0(\out[1508]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[825] ),
        .I2(\out[1572]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[399] ),
        .I4(\out[1508]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1508]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1508]_i_2 
       (.I0(\f_permutation_l_/round_in [1208]),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1592]),
        .I4(\out[1572]_i_6_n_0 ),
        .O(\out[1508]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1508]_i_3 
       (.I0(\out[1596]_i_7_n_0 ),
        .I1(padder_out_1[439]),
        .I2(out[375]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1550]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1294]),
        .O(\out[1508]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1509]_i_1 
       (.I0(\out[1509]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[826] ),
        .I2(\out[1573]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[400] ),
        .I4(\out[1509]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1509]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1509]_i_2 
       (.I0(\f_permutation_l_/round_in [1209]),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1593]),
        .I4(\out[1573]_i_6_n_0 ),
        .O(\out[1509]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1509]_i_3 
       (.I0(\out[1597]_i_7_n_0 ),
        .I1(padder_out_1[424]),
        .I2(out[360]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1551]_i_15_n_0 ),
        .I5(\f_permutation_l_/round_in [1295]),
        .O(\out[1509]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[150]_i_1 
       (.I0(\out[1469]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[687] ),
        .I2(\out[150]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[212] ),
        .I4(\out[1280]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [150]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[150]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[621] ),
        .I1(\f_permutation_l_/round_in [1516]),
        .I2(\out[1559]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[150]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[1510]_i_1 
       (.I0(\out[1510]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[827] ),
        .I2(\out[1574]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[401] ),
        .I4(\out[1510]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1510]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1510]_i_2 
       (.I0(\f_permutation_l_/round_in [1210]),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1594]),
        .I4(\out[1574]_i_6_n_0 ),
        .O(\out[1510]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1510]_i_3 
       (.I0(\out[1598]_i_7_n_0 ),
        .I1(padder_out_1[425]),
        .I2(out[361]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1552]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1296]),
        .O(\out[1510]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[1511]_i_1 
       (.I0(\out[1511]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[828] ),
        .I2(\out[1575]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[402] ),
        .I4(\out[1511]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1511]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1511]_i_2 
       (.I0(\f_permutation_l_/round_in [1211]),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1595]),
        .I4(\out[1575]_i_6_n_0 ),
        .O(\out[1511]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1511]_i_3 
       (.I0(\out[1543]_i_12_n_0 ),
        .I1(out[362]),
        .I2(padder_out_1[426]),
        .I3(\out[1599]_i_7_n_0 ),
        .I4(\out[1553]_i_14_n_0 ),
        .I5(\f_permutation_l_/round_in [1297]),
        .O(\out[1511]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[1512]_i_1 
       (.I0(\out[1512]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[829] ),
        .I2(\out[1576]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[403] ),
        .I4(\out[1512]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1512]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1512]_i_2 
       (.I0(\f_permutation_l_/round_in [1212]),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1596]),
        .I4(\out[1576]_i_6_n_0 ),
        .O(\out[1512]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1512]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[234]),
        .I2(padder_out_1[298]),
        .I3(\out[1554]_i_14_n_0 ),
        .I4(\out[1536]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1427]),
        .O(\out[1512]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[1513]_i_1 
       (.I0(\out[1513]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[830] ),
        .I2(\out[1577]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[404] ),
        .I4(\out[1513]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1513]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1513]_i_2 
       (.I0(\f_permutation_l_/round_in [1213]),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1597]),
        .I4(\out[1577]_i_6_n_0 ),
        .O(\out[1513]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1513]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[235]),
        .I2(padder_out_1[299]),
        .I3(\out[1555]_i_14_n_0 ),
        .I4(\out[1537]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1428]),
        .O(\out[1513]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[1514]_i_1 
       (.I0(\out[1514]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[831] ),
        .I2(\out[1578]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[405] ),
        .I4(\out[1514]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1514]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1514]_i_2 
       (.I0(\f_permutation_l_/round_in [1214]),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1598]),
        .I4(\out[1578]_i_6_n_0 ),
        .O(\out[1514]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1514]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[236]),
        .I2(padder_out_1[300]),
        .I3(\out[1556]_i_14_n_0 ),
        .I4(\out[1538]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1429]),
        .O(\out[1514]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[1515]_i_1 
       (.I0(\out[1515]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[768] ),
        .I2(\out[1579]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[406] ),
        .I4(\out[1515]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1515]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1515]_i_2 
       (.I0(\f_permutation_l_/round_in [1215]),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1599]),
        .I4(\out[1579]_i_7_n_0 ),
        .O(\out[1515]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h936C6C936C93936C)) 
    \out[1515]_i_3 
       (.I0(\out[1542]_i_8_n_0 ),
        .I1(out[237]),
        .I2(padder_out_1[301]),
        .I3(\out[1557]_i_13_n_0 ),
        .I4(\out[1539]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1430]),
        .O(\out[1515]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1516]_i_1 
       (.I0(\out[1516]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[769] ),
        .I2(\out[1580]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[407] ),
        .I4(\out[1516]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1516]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1516]_i_2 
       (.I0(\f_permutation_l_/round_in [1152]),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1536]),
        .I4(\out[1580]_i_6_n_0 ),
        .O(\out[1516]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1516]_i_3 
       (.I0(\out[1558]_i_14_n_0 ),
        .I1(padder_out_1[302]),
        .I2(out[238]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1540]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1431]),
        .O(\out[1516]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1517]_i_1 
       (.I0(\out[1517]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[770] ),
        .I2(\out[1581]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[408] ),
        .I4(\out[1517]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1517]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1517]_i_2 
       (.I0(\f_permutation_l_/round_in [1153]),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1537]),
        .I4(\out[1581]_i_6_n_0 ),
        .O(\out[1517]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1517]_i_3 
       (.I0(\out[1559]_i_15_n_0 ),
        .I1(padder_out_1[303]),
        .I2(out[239]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1541]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1432]),
        .O(\out[1517]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1518]_i_1 
       (.I0(\out[1518]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[771] ),
        .I2(\out[1582]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[409] ),
        .I4(\out[1518]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1518]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1518]_i_2 
       (.I0(\f_permutation_l_/round_in [1154]),
        .I1(\f_permutation_l_/round_in [1409]),
        .I2(\out[1582]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1538]),
        .I4(\out[1582]_i_6_n_0 ),
        .O(\out[1518]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1518]_i_3 
       (.I0(\out[1560]_i_15_n_0 ),
        .I1(padder_out_1[288]),
        .I2(out[224]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1542]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1433]),
        .O(\out[1518]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1519]_i_1 
       (.I0(\out[1519]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[772] ),
        .I2(\out[1583]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[410] ),
        .I4(\out[1519]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1519]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1519]_i_2 
       (.I0(\f_permutation_l_/round_in [1155]),
        .I1(\f_permutation_l_/round_in [1410]),
        .I2(\out[1583]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1539]),
        .I4(\out[1583]_i_6_n_0 ),
        .O(\out[1519]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1519]_i_3 
       (.I0(\out[1561]_i_14_n_0 ),
        .I1(padder_out_1[289]),
        .I2(out[225]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1543]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1434]),
        .O(\out[1519]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[151]_i_1 
       (.I0(\out[1470]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[688] ),
        .I2(\out[151]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[213] ),
        .I4(\out[1281]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [151]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[151]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[622] ),
        .I1(\f_permutation_l_/round_in [1517]),
        .I2(\out[1560]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[151]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1520]_i_1 
       (.I0(\out[1520]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[773] ),
        .I2(\out[1584]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[411] ),
        .I4(\out[1520]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1520]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1520]_i_2 
       (.I0(\f_permutation_l_/round_in [1156]),
        .I1(\f_permutation_l_/round_in [1411]),
        .I2(\out[1584]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1540]),
        .I4(\out[1584]_i_6_n_0 ),
        .O(\out[1520]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1520]_i_3 
       (.I0(\out[1562]_i_15_n_0 ),
        .I1(padder_out_1[290]),
        .I2(out[226]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1544]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1435]),
        .O(\out[1520]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1521]_i_1 
       (.I0(\out[1521]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[774] ),
        .I2(\out[1585]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[412] ),
        .I4(\out[1521]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1521]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1521]_i_2 
       (.I0(\f_permutation_l_/round_in [1157]),
        .I1(\f_permutation_l_/round_in [1412]),
        .I2(\out[1585]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1541]),
        .I4(\out[1585]_i_6_n_0 ),
        .O(\out[1521]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1521]_i_3 
       (.I0(\out[1563]_i_14_n_0 ),
        .I1(padder_out_1[291]),
        .I2(out[227]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1545]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1436]),
        .O(\out[1521]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1522]_i_1 
       (.I0(\out[1522]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[775] ),
        .I2(\out[1586]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[413] ),
        .I4(\out[1522]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1522]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1522]_i_2 
       (.I0(\f_permutation_l_/round_in [1158]),
        .I1(\f_permutation_l_/round_in [1413]),
        .I2(\out[1586]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1542]),
        .I4(\out[1586]_i_6_n_0 ),
        .O(\out[1522]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1522]_i_3 
       (.I0(\out[1564]_i_15_n_0 ),
        .I1(padder_out_1[292]),
        .I2(out[228]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1546]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1437]),
        .O(\out[1522]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1523]_i_1 
       (.I0(\out[1523]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[776] ),
        .I2(\out[1587]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[414] ),
        .I4(\out[1523]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1523]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1523]_i_2 
       (.I0(\f_permutation_l_/round_in [1159]),
        .I1(\f_permutation_l_/round_in [1414]),
        .I2(\out[1587]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1543]),
        .I4(\out[1587]_i_6_n_0 ),
        .O(\out[1523]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1523]_i_3 
       (.I0(\out[1565]_i_15_n_0 ),
        .I1(padder_out_1[293]),
        .I2(out[229]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1547]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1438]),
        .O(\out[1523]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1524]_i_1 
       (.I0(\out[1524]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[777] ),
        .I2(\out[1588]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[415] ),
        .I4(\out[1524]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1524]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1524]_i_2 
       (.I0(\f_permutation_l_/round_in [1160]),
        .I1(\f_permutation_l_/round_in [1415]),
        .I2(\out[1588]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1544]),
        .I4(\out[1588]_i_6_n_0 ),
        .O(\out[1524]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1524]_i_3 
       (.I0(\out[1566]_i_14_n_0 ),
        .I1(padder_out_1[294]),
        .I2(out[230]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1548]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1439]),
        .O(\out[1524]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1525]_i_1 
       (.I0(\out[1525]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[778] ),
        .I2(\out[1589]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[416] ),
        .I4(\out[1525]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1525]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1525]_i_2 
       (.I0(\f_permutation_l_/round_in [1161]),
        .I1(\f_permutation_l_/round_in [1416]),
        .I2(\out[1589]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1545]),
        .I4(\out[1589]_i_6_n_0 ),
        .O(\out[1525]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1525]_i_3 
       (.I0(\out[1567]_i_16_n_0 ),
        .I1(padder_out_1[295]),
        .I2(out[231]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1549]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1440]),
        .O(\out[1525]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1526]_i_1 
       (.I0(\out[1526]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[779] ),
        .I2(\out[1590]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[417] ),
        .I4(\out[1526]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1526]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1526]_i_2 
       (.I0(\f_permutation_l_/round_in [1162]),
        .I1(\f_permutation_l_/round_in [1417]),
        .I2(\out[1590]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1546]),
        .I4(\out[1590]_i_6_n_0 ),
        .O(\out[1526]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1526]_i_3 
       (.I0(\out[1568]_i_15_n_0 ),
        .I1(padder_out_1[280]),
        .I2(out[216]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1550]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1441]),
        .O(\out[1526]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1527]_i_1 
       (.I0(\out[1527]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[780] ),
        .I2(\out[1591]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[418] ),
        .I4(\out[1527]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1527]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1527]_i_2 
       (.I0(\f_permutation_l_/round_in [1163]),
        .I1(\f_permutation_l_/round_in [1418]),
        .I2(\out[1591]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1547]),
        .I4(\out[1591]_i_6_n_0 ),
        .O(\out[1527]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1527]_i_3 
       (.I0(\out[1569]_i_15_n_0 ),
        .I1(padder_out_1[281]),
        .I2(out[217]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1551]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1442]),
        .O(\out[1527]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1528]_i_1 
       (.I0(\out[1528]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[781] ),
        .I2(\out[1592]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[419] ),
        .I4(\out[1528]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1528]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1528]_i_2 
       (.I0(\f_permutation_l_/round_in [1164]),
        .I1(\f_permutation_l_/round_in [1419]),
        .I2(\out[1592]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1548]),
        .I4(\out[1592]_i_6_n_0 ),
        .O(\out[1528]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1528]_i_3 
       (.I0(\out[1570]_i_15_n_0 ),
        .I1(padder_out_1[282]),
        .I2(out[218]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1552]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1443]),
        .O(\out[1528]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1529]_i_1 
       (.I0(\out[1529]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[782] ),
        .I2(\out[1593]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[420] ),
        .I4(\out[1529]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1529]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1529]_i_2 
       (.I0(\f_permutation_l_/round_in [1165]),
        .I1(\f_permutation_l_/round_in [1420]),
        .I2(\out[1593]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1549]),
        .I4(\out[1593]_i_6_n_0 ),
        .O(\out[1529]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1529]_i_3 
       (.I0(\out[1571]_i_14_n_0 ),
        .I1(padder_out_1[283]),
        .I2(out[219]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1553]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1444]),
        .O(\out[1529]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[152]_i_1 
       (.I0(\out[1471]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[689] ),
        .I2(\out[152]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[214] ),
        .I4(\out[1538]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [152]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[152]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[623] ),
        .I1(\f_permutation_l_/round_in [1518]),
        .I2(\out[1561]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[152]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1530]_i_1 
       (.I0(\out[1530]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[783] ),
        .I2(\out[1594]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[421] ),
        .I4(\out[1530]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1530]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1530]_i_2 
       (.I0(\f_permutation_l_/round_in [1166]),
        .I1(\f_permutation_l_/round_in [1421]),
        .I2(\out[1594]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1550]),
        .I4(\out[1594]_i_6_n_0 ),
        .O(\out[1530]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1530]_i_3 
       (.I0(\out[1572]_i_15_n_0 ),
        .I1(padder_out_1[284]),
        .I2(out[220]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1554]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1445]),
        .O(\out[1530]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1531]_i_1 
       (.I0(\out[1531]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[784] ),
        .I2(\out[1595]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[422] ),
        .I4(\out[1531]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1531]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1531]_i_2 
       (.I0(\f_permutation_l_/round_in [1167]),
        .I1(\f_permutation_l_/round_in [1422]),
        .I2(\out[1595]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1551]),
        .I4(\out[1595]_i_6_n_0 ),
        .O(\out[1531]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1531]_i_3 
       (.I0(\out[1573]_i_15_n_0 ),
        .I1(padder_out_1[285]),
        .I2(out[221]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1555]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1446]),
        .O(\out[1531]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1532]_i_1 
       (.I0(\out[1532]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[785] ),
        .I2(\out[1596]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[423] ),
        .I4(\out[1532]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1532]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1532]_i_2 
       (.I0(\f_permutation_l_/round_in [1168]),
        .I1(\f_permutation_l_/round_in [1423]),
        .I2(\out[1596]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1552]),
        .I4(\out[1596]_i_6_n_0 ),
        .O(\out[1532]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1532]_i_3 
       (.I0(\out[1574]_i_15_n_0 ),
        .I1(padder_out_1[286]),
        .I2(out[222]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1556]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1447]),
        .O(\out[1532]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1533]_i_1 
       (.I0(\out[1533]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[786] ),
        .I2(\out[1597]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[424] ),
        .I4(\out[1533]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1533]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1533]_i_2 
       (.I0(\f_permutation_l_/round_in [1169]),
        .I1(\f_permutation_l_/round_in [1424]),
        .I2(\out[1597]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1553]),
        .I4(\out[1597]_i_6_n_0 ),
        .O(\out[1533]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1533]_i_3 
       (.I0(\out[1575]_i_15_n_0 ),
        .I1(padder_out_1[287]),
        .I2(out[223]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1557]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1448]),
        .O(\out[1533]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1534]_i_1 
       (.I0(\out[1534]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[787] ),
        .I2(\out[1598]_i_4_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[425] ),
        .I4(\out[1534]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [1534]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1534]_i_2 
       (.I0(\f_permutation_l_/round_in [1170]),
        .I1(\f_permutation_l_/round_in [1425]),
        .I2(\out[1598]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1554]),
        .I4(\out[1598]_i_6_n_0 ),
        .O(\out[1534]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1534]_i_3 
       (.I0(\out[1576]_i_15_n_0 ),
        .I1(padder_out_1[272]),
        .I2(out[208]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1558]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1449]),
        .O(\out[1534]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[1535]_i_1 
       (.I0(\out[1599]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[788] ),
        .I2(\out[1599]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[426] ),
        .I4(\out[1535]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1535]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1535]_i_2 
       (.I0(\out[1577]_i_15_n_0 ),
        .I1(padder_out_1[273]),
        .I2(out[209]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1559]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1450]),
        .O(\out[1535]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4B4B4B4B4B4B4BB4)) 
    \out[1536]_i_1 
       (.I0(\out[1536]_i_2_n_0 ),
        .I1(\out[1536]_i_3_n_0 ),
        .I2(\out[1536]_i_4_n_0 ),
        .I3(\out[1536]_i_5_n_0 ),
        .I4(\out[1536]_i_6_n_0 ),
        .I5(\f_permutation_l_/i_reg_n_0_[12] ),
        .O(\f_permutation_l_/round_out [1536]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1536]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[916] ),
        .I1(padder_out_1[236]),
        .I2(out[172]),
        .I3(\f_permutation_l_/out_reg_n_0_[276] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[596] ),
        .O(\out[1536]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_11 
       (.I0(padder_out_1[364]),
        .I1(out[300]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1364]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1536]_i_12 
       (.I0(\f_permutation_l_/out_reg_n_0_[724] ),
        .I1(padder_out_1[44]),
        .I2(\f_permutation_l_/out_reg_n_0_[1044] ),
        .I3(\f_permutation_l_/out_reg_n_0_[84] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[404] ),
        .O(\out[1536]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_13 
       (.I0(padder_out_1[493]),
        .I1(out[429]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1493]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1536]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[853] ),
        .I1(padder_out_1[173]),
        .I2(out[109]),
        .I3(\f_permutation_l_/out_reg_n_0_[213] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[533] ),
        .O(\out[1536]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_15 
       (.I0(padder_out_1[568]),
        .I1(out[504]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1536]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_16 
       (.I0(padder_out_1[312]),
        .I1(out[248]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1280]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1536]_i_17 
       (.I0(\f_permutation_l_/out_reg_n_0_[640] ),
        .I1(\f_permutation_l_/out_reg_n_0_[960] ),
        .I2(\f_permutation_l_/out_reg_n_0_ ),
        .I3(\f_permutation_l_/out_reg_n_0_[320] ),
        .O(\out[1536]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_18 
       (.I0(padder_out_1[455]),
        .I1(out[391]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1535]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1536]_i_19 
       (.I0(\f_permutation_l_/out_reg_n_0_[895] ),
        .I1(padder_out_1[135]),
        .I2(out[71]),
        .I3(\f_permutation_l_/out_reg_n_0_[255] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[575] ),
        .O(\out[1536]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1536]_i_2 
       (.I0(\f_permutation_l_/round_in [1172]),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1556]),
        .I4(\out[1536]_i_10_n_0 ),
        .O(\out[1536]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1536]_i_3 
       (.I0(\f_permutation_l_/out_reg_n_0_[789] ),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1493]),
        .I4(\out[1536]_i_14_n_0 ),
        .O(\out[1536]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1536]_i_4 
       (.I0(\f_permutation_l_/round_in [1536]),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[1536]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1536]_i_5 
       (.I0(\f_permutation_l_/i_reg_n_0_[21] ),
        .I1(\f_permutation_l_/i_reg_n_0_[4] ),
        .I2(update__0_i_1_n_0),
        .I3(\f_permutation_l_/i_reg_n_0_[19] ),
        .I4(\f_permutation_l_/i_reg_n_0_[5] ),
        .I5(\f_permutation_l_/i_reg_n_0_[14] ),
        .O(\out[1536]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \out[1536]_i_6 
       (.I0(\f_permutation_l_/i_reg_n_0_[9] ),
        .I1(\f_permutation_l_/i_reg_n_0_[3] ),
        .I2(\f_permutation_l_/i_reg_n_0_[11] ),
        .I3(\f_permutation_l_/i_reg_n_0_[13] ),
        .I4(\f_permutation_l_/i_reg_n_0_[6] ),
        .O(\out[1536]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_7 
       (.I0(padder_out_1[427]),
        .I1(out[363]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1427]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1536]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[787] ),
        .I1(padder_out_1[107]),
        .I2(out[43]),
        .I3(\f_permutation_l_/out_reg_n_0_[147] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[467] ),
        .O(\out[1536]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1536]_i_9 
       (.I0(padder_out_1[556]),
        .I1(out[492]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1556]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41BEBE41)) 
    \out[1537]_i_1 
       (.I0(\out[1537]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[790] ),
        .I2(\out[1537]_i_3_n_0 ),
        .I3(\out[1537]_i_4_n_0 ),
        .I4(\f_permutation_l_/rc [1]),
        .O(\f_permutation_l_/round_out [1537]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1537]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[854] ),
        .I1(padder_out_1[174]),
        .I2(out[110]),
        .I3(\f_permutation_l_/out_reg_n_0_[214] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[534] ),
        .O(\out[1537]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1537]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[725] ),
        .I1(padder_out_1[45]),
        .I2(\f_permutation_l_/out_reg_n_0_[1045] ),
        .I3(\f_permutation_l_/out_reg_n_0_[85] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[405] ),
        .O(\out[1537]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_12 
       (.I0(padder_out_1[365]),
        .I1(out[301]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1365]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_13 
       (.I0(padder_out_1[569]),
        .I1(out[505]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1537]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_14 
       (.I0(padder_out_1[313]),
        .I1(out[249]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1281]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1537]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[641] ),
        .I1(\f_permutation_l_/out_reg_n_0_[961] ),
        .I2(\f_permutation_l_/out_reg_n_0_[1] ),
        .I3(\f_permutation_l_/out_reg_n_0_[321] ),
        .O(\out[1537]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_16 
       (.I0(padder_out_1[504]),
        .I1(out[440]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1472]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1537]_i_17 
       (.I0(\f_permutation_l_/out_reg_n_0_[832] ),
        .I1(padder_out_1[184]),
        .I2(out[120]),
        .I3(\f_permutation_l_/out_reg_n_0_[192] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[512] ),
        .O(\out[1537]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \out[1537]_i_18 
       (.I0(\f_permutation_l_/i_reg_n_0_[14] ),
        .I1(\f_permutation_l_/i_reg_n_0_[15] ),
        .O(\out[1537]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1537]_i_2 
       (.I0(\f_permutation_l_/round_in [1173]),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1557]),
        .I4(\out[1537]_i_9_n_0 ),
        .O(\out[1537]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1537]_i_3 
       (.I0(\out[1537]_i_10_n_0 ),
        .I1(padder_out_1[494]),
        .I2(out[430]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1537]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1365]),
        .O(\out[1537]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1537]_i_4 
       (.I0(\f_permutation_l_/round_in [1537]),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[1537]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1537]_i_5 
       (.I0(\out[1543]_i_22_n_0 ),
        .I1(\f_permutation_l_/i_reg_n_0_[18] ),
        .I2(\f_permutation_l_/i_reg_n_0_[10] ),
        .I3(\out[1537]_i_18_n_0 ),
        .I4(\f_permutation_l_/i_reg_n_0_[17] ),
        .I5(\out[1543]_i_20_n_0 ),
        .O(\f_permutation_l_/rc [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_6 
       (.I0(padder_out_1[428]),
        .I1(out[364]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1428]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1537]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[788] ),
        .I1(padder_out_1[108]),
        .I2(out[44]),
        .I3(\f_permutation_l_/out_reg_n_0_[148] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[468] ),
        .O(\out[1537]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1537]_i_8 
       (.I0(padder_out_1[557]),
        .I1(out[493]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1557]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1537]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[917] ),
        .I1(padder_out_1[237]),
        .I2(out[173]),
        .I3(\f_permutation_l_/out_reg_n_0_[277] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[597] ),
        .O(\out[1537]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1538]_i_1 
       (.I0(\f_permutation_l_/round_in [1174]),
        .I1(\out[1538]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[791] ),
        .I3(\out[1538]_i_4_n_0 ),
        .I4(\out[1538]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1538]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1538]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[726] ),
        .I1(padder_out_1[46]),
        .I2(\f_permutation_l_/out_reg_n_0_[1046] ),
        .I3(\f_permutation_l_/out_reg_n_0_[86] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[406] ),
        .O(\out[1538]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_11 
       (.I0(padder_out_1[366]),
        .I1(out[302]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1366]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_12 
       (.I0(padder_out_1[570]),
        .I1(out[506]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1538]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_13 
       (.I0(padder_out_1[314]),
        .I1(out[250]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1282]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1538]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[642] ),
        .I1(\f_permutation_l_/out_reg_n_0_[962] ),
        .I2(\f_permutation_l_/out_reg_n_0_[2] ),
        .I3(\f_permutation_l_/out_reg_n_0_[322] ),
        .O(\out[1538]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_15 
       (.I0(padder_out_1[505]),
        .I1(out[441]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1473]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1538]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[833] ),
        .I1(padder_out_1[185]),
        .I2(out[121]),
        .I3(\f_permutation_l_/out_reg_n_0_[193] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[513] ),
        .O(\out[1538]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_2 
       (.I0(padder_out_1[174]),
        .I1(out[110]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1174]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1538]_i_3 
       (.I0(\out[1538]_i_6_n_0 ),
        .I1(padder_out_1[558]),
        .I2(out[494]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1538]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1429]),
        .O(\out[1538]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1538]_i_4 
       (.I0(\out[1538]_i_9_n_0 ),
        .I1(padder_out_1[495]),
        .I2(out[431]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1538]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1366]),
        .O(\out[1538]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1538]_i_5 
       (.I0(\f_permutation_l_/round_in [1538]),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[1538]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1538]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[918] ),
        .I1(padder_out_1[238]),
        .I2(out[174]),
        .I3(\f_permutation_l_/out_reg_n_0_[278] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[598] ),
        .O(\out[1538]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1538]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[789] ),
        .I1(padder_out_1[109]),
        .I2(out[45]),
        .I3(\f_permutation_l_/out_reg_n_0_[149] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[469] ),
        .O(\out[1538]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1538]_i_8 
       (.I0(padder_out_1[429]),
        .I1(out[365]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1429]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1538]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[855] ),
        .I1(padder_out_1[175]),
        .I2(out[111]),
        .I3(\f_permutation_l_/out_reg_n_0_[215] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[535] ),
        .O(\out[1538]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h906F6F906F90906F)) 
    \out[1539]_i_1 
       (.I0(\f_permutation_l_/round_in [1175]),
        .I1(\out[1539]_i_3_n_0 ),
        .I2(\out[1539]_i_4_n_0 ),
        .I3(\f_permutation_l_/round_in [1539]),
        .I4(\out[1539]_i_6_n_0 ),
        .I5(\f_permutation_l_/rc [3]),
        .O(\f_permutation_l_/round_out [1539]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_10 
       (.I0(padder_out_1[430]),
        .I1(out[366]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1430]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_11 
       (.I0(padder_out_1[367]),
        .I1(out[303]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1367]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1539]_i_12 
       (.I0(\f_permutation_l_/out_reg_n_0_[727] ),
        .I1(padder_out_1[47]),
        .I2(\f_permutation_l_/out_reg_n_0_[1047] ),
        .I3(\f_permutation_l_/out_reg_n_0_[87] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[407] ),
        .O(\out[1539]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_13 
       (.I0(padder_out_1[480]),
        .I1(out[416]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1496]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1539]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[856] ),
        .I1(padder_out_1[160]),
        .I2(out[96]),
        .I3(\f_permutation_l_/out_reg_n_0_[216] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[536] ),
        .O(\out[1539]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1539]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[834] ),
        .I1(padder_out_1[186]),
        .I2(out[122]),
        .I3(\f_permutation_l_/out_reg_n_0_[194] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[514] ),
        .O(\out[1539]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1539]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[643] ),
        .I1(\f_permutation_l_/out_reg_n_0_[963] ),
        .I2(\f_permutation_l_/out_reg_n_0_[3] ),
        .I3(\f_permutation_l_/out_reg_n_0_[323] ),
        .O(\out[1539]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_17 
       (.I0(padder_out_1[315]),
        .I1(out[251]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1283]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \out[1539]_i_18 
       (.I0(\f_permutation_l_/i_reg_n_0_[10] ),
        .I1(\f_permutation_l_/i_reg_n_0_[18] ),
        .O(\out[1539]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_2 
       (.I0(padder_out_1[175]),
        .I1(out[111]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1175]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1539]_i_3 
       (.I0(\out[1539]_i_8_n_0 ),
        .I1(padder_out_1[559]),
        .I2(out[495]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1539]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1430]),
        .O(\out[1539]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1539]_i_4 
       (.I0(\f_permutation_l_/out_reg_n_0_[792] ),
        .I1(\f_permutation_l_/round_in [1367]),
        .I2(\out[1539]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1496]),
        .I4(\out[1539]_i_14_n_0 ),
        .O(\out[1539]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1539]_i_5 
       (.I0(padder_out_1[571]),
        .I1(out[507]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1539]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1539]_i_6 
       (.I0(\out[1539]_i_15_n_0 ),
        .I1(padder_out_1[506]),
        .I2(out[442]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1539]_i_16_n_0 ),
        .I5(\f_permutation_l_/round_in [1283]),
        .O(\out[1539]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1539]_i_7 
       (.I0(\out[1543]_i_20_n_0 ),
        .I1(\f_permutation_l_/i_reg_n_0_[17] ),
        .I2(\f_permutation_l_/i_reg_n_0_[8] ),
        .I3(\out[1539]_i_18_n_0 ),
        .I4(\out[1536]_i_6_n_0 ),
        .I5(\f_permutation_l_/p_0_in ),
        .O(\f_permutation_l_/rc [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1539]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[919] ),
        .I1(padder_out_1[239]),
        .I2(out[175]),
        .I3(\f_permutation_l_/out_reg_n_0_[279] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[599] ),
        .O(\out[1539]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1539]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[790] ),
        .I1(padder_out_1[110]),
        .I2(out[46]),
        .I3(\f_permutation_l_/out_reg_n_0_[150] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[470] ),
        .O(\out[1539]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[153]_i_1 
       (.I0(\out[1408]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[690] ),
        .I2(\out[153]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[215] ),
        .I4(\out[1539]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [153]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[153]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[624] ),
        .I1(\f_permutation_l_/round_in [1519]),
        .I2(\out[1562]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[153]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1540]_i_1 
       (.I0(\f_permutation_l_/round_in [1176]),
        .I1(\out[1540]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[793] ),
        .I3(\out[1540]_i_4_n_0 ),
        .I4(\out[1540]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1540]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1540]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[728] ),
        .I1(padder_out_1[32]),
        .I2(\f_permutation_l_/out_reg_n_0_[1048] ),
        .I3(\f_permutation_l_/out_reg_n_0_[88] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[408] ),
        .O(\out[1540]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_11 
       (.I0(padder_out_1[352]),
        .I1(out[288]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1368]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_12 
       (.I0(padder_out_1[572]),
        .I1(out[508]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1540]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_13 
       (.I0(padder_out_1[316]),
        .I1(out[252]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1284]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1540]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[644] ),
        .I1(\f_permutation_l_/out_reg_n_0_[964] ),
        .I2(\f_permutation_l_/out_reg_n_0_[4] ),
        .I3(\f_permutation_l_/out_reg_n_0_[324] ),
        .O(\out[1540]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_15 
       (.I0(padder_out_1[507]),
        .I1(out[443]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1475]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1540]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[835] ),
        .I1(padder_out_1[187]),
        .I2(out[123]),
        .I3(\f_permutation_l_/out_reg_n_0_[195] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[515] ),
        .O(\out[1540]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_2 
       (.I0(padder_out_1[160]),
        .I1(out[96]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1176]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1540]_i_3 
       (.I0(\out[1540]_i_6_n_0 ),
        .I1(padder_out_1[544]),
        .I2(out[480]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1540]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1431]),
        .O(\out[1540]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1540]_i_4 
       (.I0(\out[1540]_i_9_n_0 ),
        .I1(padder_out_1[481]),
        .I2(out[417]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1540]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1368]),
        .O(\out[1540]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1540]_i_5 
       (.I0(\f_permutation_l_/round_in [1540]),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[1540]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1540]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[920] ),
        .I1(padder_out_1[224]),
        .I2(out[160]),
        .I3(\f_permutation_l_/out_reg_n_0_[280] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[600] ),
        .O(\out[1540]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1540]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[791] ),
        .I1(padder_out_1[111]),
        .I2(out[47]),
        .I3(\f_permutation_l_/out_reg_n_0_[151] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[471] ),
        .O(\out[1540]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1540]_i_8 
       (.I0(padder_out_1[431]),
        .I1(out[367]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1431]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1540]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[857] ),
        .I1(padder_out_1[161]),
        .I2(out[97]),
        .I3(\f_permutation_l_/out_reg_n_0_[217] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[537] ),
        .O(\out[1540]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1541]_i_1 
       (.I0(\f_permutation_l_/round_in [1177]),
        .I1(\out[1541]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[794] ),
        .I3(\out[1541]_i_4_n_0 ),
        .I4(\out[1541]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1541]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1541]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[729] ),
        .I1(padder_out_1[33]),
        .I2(\f_permutation_l_/out_reg_n_0_[1049] ),
        .I3(\f_permutation_l_/out_reg_n_0_[89] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[409] ),
        .O(\out[1541]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_11 
       (.I0(padder_out_1[353]),
        .I1(out[289]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1369]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_12 
       (.I0(padder_out_1[573]),
        .I1(out[509]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1541]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_13 
       (.I0(padder_out_1[317]),
        .I1(out[253]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1285]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1541]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[645] ),
        .I1(\f_permutation_l_/out_reg_n_0_[965] ),
        .I2(\f_permutation_l_/out_reg_n_0_[5] ),
        .I3(\f_permutation_l_/out_reg_n_0_[325] ),
        .O(\out[1541]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_15 
       (.I0(padder_out_1[508]),
        .I1(out[444]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1476]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1541]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[836] ),
        .I1(padder_out_1[188]),
        .I2(out[124]),
        .I3(\f_permutation_l_/out_reg_n_0_[196] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[516] ),
        .O(\out[1541]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_2 
       (.I0(padder_out_1[161]),
        .I1(out[97]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1177]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1541]_i_3 
       (.I0(\out[1541]_i_6_n_0 ),
        .I1(padder_out_1[545]),
        .I2(out[481]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1541]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1432]),
        .O(\out[1541]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1541]_i_4 
       (.I0(\out[1541]_i_9_n_0 ),
        .I1(padder_out_1[482]),
        .I2(out[418]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1541]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1369]),
        .O(\out[1541]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1541]_i_5 
       (.I0(\f_permutation_l_/round_in [1541]),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[1541]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1541]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[921] ),
        .I1(padder_out_1[225]),
        .I2(out[161]),
        .I3(\f_permutation_l_/out_reg_n_0_[281] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[601] ),
        .O(\out[1541]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1541]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[792] ),
        .I1(padder_out_1[96]),
        .I2(out[32]),
        .I3(\f_permutation_l_/out_reg_n_0_[152] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[472] ),
        .O(\out[1541]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1541]_i_8 
       (.I0(padder_out_1[416]),
        .I1(out[352]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1432]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1541]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[858] ),
        .I1(padder_out_1[162]),
        .I2(out[98]),
        .I3(\f_permutation_l_/out_reg_n_0_[218] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[538] ),
        .O(\out[1541]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1542]_i_1 
       (.I0(\f_permutation_l_/round_in [1178]),
        .I1(\out[1542]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[795] ),
        .I3(\out[1542]_i_4_n_0 ),
        .I4(\out[1542]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1542]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_10 
       (.I0(padder_out_1[417]),
        .I1(out[353]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1433]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1542]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[859] ),
        .I1(padder_out_1[163]),
        .I2(out[99]),
        .I3(\f_permutation_l_/out_reg_n_0_[219] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[539] ),
        .O(\out[1542]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1542]_i_12 
       (.I0(\f_permutation_l_/out_reg_n_0_[730] ),
        .I1(padder_out_1[34]),
        .I2(\f_permutation_l_/out_reg_n_0_[1050] ),
        .I3(\f_permutation_l_/out_reg_n_0_[90] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[410] ),
        .O(\out[1542]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_13 
       (.I0(padder_out_1[354]),
        .I1(out[290]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1370]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_14 
       (.I0(padder_out_1[574]),
        .I1(out[510]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1542]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_15 
       (.I0(padder_out_1[318]),
        .I1(out[254]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1286]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1542]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[646] ),
        .I1(\f_permutation_l_/out_reg_n_0_[966] ),
        .I2(\f_permutation_l_/out_reg_n_0_[6] ),
        .I3(\f_permutation_l_/out_reg_n_0_[326] ),
        .O(\out[1542]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_17 
       (.I0(padder_out_1[509]),
        .I1(out[445]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1477]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1542]_i_18 
       (.I0(\f_permutation_l_/out_reg_n_0_[837] ),
        .I1(padder_out_1[189]),
        .I2(out[125]),
        .I3(\f_permutation_l_/out_reg_n_0_[197] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[517] ),
        .O(\out[1542]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1542]_i_2 
       (.I0(padder_out_1[162]),
        .I1(out[98]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1178]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1542]_i_3 
       (.I0(\out[1542]_i_7_n_0 ),
        .I1(padder_out_1[546]),
        .I2(out[482]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1542]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1433]),
        .O(\out[1542]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1542]_i_4 
       (.I0(\out[1542]_i_11_n_0 ),
        .I1(padder_out_1[483]),
        .I2(out[419]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1542]_i_12_n_0 ),
        .I5(\f_permutation_l_/round_in [1370]),
        .O(\out[1542]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1542]_i_5 
       (.I0(\f_permutation_l_/round_in [1542]),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[1542]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1542]_i_6 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1542]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1542]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[922] ),
        .I1(padder_out_1[226]),
        .I2(out[162]),
        .I3(\f_permutation_l_/out_reg_n_0_[282] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[602] ),
        .O(\out[1542]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1542]_i_8 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1542]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1542]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[793] ),
        .I1(padder_out_1[97]),
        .I2(out[33]),
        .I3(\f_permutation_l_/out_reg_n_0_[153] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[473] ),
        .O(\out[1542]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \out[1543]_i_1 
       (.I0(\f_permutation_l_/calc ),
        .I1(update__0_i_1_n_0),
        .O(\f_permutation_l_/update ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1543]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[923] ),
        .I1(padder_out_1[227]),
        .I2(out[163]),
        .I3(\f_permutation_l_/out_reg_n_0_[283] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[603] ),
        .O(\out[1543]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1543]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[860] ),
        .I1(padder_out_1[164]),
        .I2(out[100]),
        .I3(\f_permutation_l_/out_reg_n_0_[220] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[540] ),
        .O(\out[1543]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1543]_i_12 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1543]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1543]_i_13 
       (.I0(\f_permutation_l_/out_reg_n_0_[731] ),
        .I1(padder_out_1[35]),
        .I2(\f_permutation_l_/out_reg_n_0_[1051] ),
        .I3(\f_permutation_l_/out_reg_n_0_[91] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[411] ),
        .O(\out[1543]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_14 
       (.I0(padder_out_1[355]),
        .I1(out[291]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1371]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_15 
       (.I0(padder_out_1[575]),
        .I1(out[511]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1543]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_16 
       (.I0(padder_out_1[319]),
        .I1(out[255]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1287]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1543]_i_17 
       (.I0(\f_permutation_l_/out_reg_n_0_[647] ),
        .I1(\f_permutation_l_/out_reg_n_0_[967] ),
        .I2(\f_permutation_l_/out_reg_n_0_[7] ),
        .I3(\f_permutation_l_/out_reg_n_0_[327] ),
        .O(\out[1543]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_18 
       (.I0(padder_out_1[510]),
        .I1(out[446]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1478]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1543]_i_19 
       (.I0(\f_permutation_l_/out_reg_n_0_[838] ),
        .I1(padder_out_1[190]),
        .I2(out[126]),
        .I3(\f_permutation_l_/out_reg_n_0_[198] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[518] ),
        .O(\out[1543]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41BEBE41)) 
    \out[1543]_i_2 
       (.I0(\out[1543]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[796] ),
        .I2(\out[1543]_i_4_n_0 ),
        .I3(\out[1543]_i_5_n_0 ),
        .I4(\f_permutation_l_/rc [7]),
        .O(\f_permutation_l_/round_out [1543]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \out[1543]_i_20 
       (.I0(\f_permutation_l_/i_reg_n_0_[12] ),
        .I1(\f_permutation_l_/i_reg_n_0_[1] ),
        .I2(\f_permutation_l_/i_reg_n_0_[7] ),
        .O(\out[1543]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \out[1543]_i_21 
       (.I0(\f_permutation_l_/i_reg_n_0_[5] ),
        .I1(\f_permutation_l_/i_reg_n_0_[19] ),
        .I2(\f_permutation_l_/i_reg_n_0_[20] ),
        .O(\out[1543]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \out[1543]_i_22 
       (.I0(\f_permutation_l_/i_reg_n_0_ ),
        .I1(\f_permutation_l_/i_reg_n_0_[11] ),
        .I2(\f_permutation_l_/i_reg_n_0_[3] ),
        .O(\out[1543]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1543]_i_23 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1543]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1543]_i_3 
       (.I0(\f_permutation_l_/round_in [1179]),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1563]),
        .I4(\out[1543]_i_10_n_0 ),
        .O(\out[1543]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1543]_i_4 
       (.I0(\out[1543]_i_11_n_0 ),
        .I1(padder_out_1[484]),
        .I2(out[420]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1543]_i_13_n_0 ),
        .I5(\f_permutation_l_/round_in [1371]),
        .O(\out[1543]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1543]_i_5 
       (.I0(\f_permutation_l_/round_in [1543]),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[1543]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1543]_i_6 
       (.I0(\f_permutation_l_/i_reg_n_0_[8] ),
        .I1(\f_permutation_l_/i_reg_n_0_[16] ),
        .I2(\f_permutation_l_/i_reg_n_0_[13] ),
        .I3(\out[1543]_i_20_n_0 ),
        .I4(\out[1543]_i_21_n_0 ),
        .I5(\out[1543]_i_22_n_0 ),
        .O(\f_permutation_l_/rc [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_7 
       (.I0(padder_out_1[418]),
        .I1(out[354]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1434]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1543]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[794] ),
        .I1(padder_out_1[98]),
        .I2(out[34]),
        .I3(\f_permutation_l_/out_reg_n_0_[154] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[474] ),
        .O(\out[1543]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1543]_i_9 
       (.I0(padder_out_1[547]),
        .I1(out[483]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1563]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1544]_i_1 
       (.I0(\f_permutation_l_/round_in [1180]),
        .I1(\out[1544]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[797] ),
        .I3(\out[1544]_i_4_n_0 ),
        .I4(\out[1544]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1544]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1544]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[732] ),
        .I1(padder_out_1[36]),
        .I2(\f_permutation_l_/out_reg_n_0_[1052] ),
        .I3(\f_permutation_l_/out_reg_n_0_[92] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[412] ),
        .O(\out[1544]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_11 
       (.I0(padder_out_1[356]),
        .I1(out[292]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1372]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_12 
       (.I0(padder_out_1[560]),
        .I1(out[496]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1544]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_13 
       (.I0(padder_out_1[304]),
        .I1(out[240]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1288]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1544]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[648] ),
        .I1(\f_permutation_l_/out_reg_n_0_[968] ),
        .I2(\f_permutation_l_/out_reg_n_0_[8] ),
        .I3(\f_permutation_l_/out_reg_n_0_[328] ),
        .O(\out[1544]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_15 
       (.I0(padder_out_1[511]),
        .I1(out[447]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1479]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1544]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[839] ),
        .I1(padder_out_1[191]),
        .I2(out[127]),
        .I3(\f_permutation_l_/out_reg_n_0_[199] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[519] ),
        .O(\out[1544]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_2 
       (.I0(padder_out_1[164]),
        .I1(out[100]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1180]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1544]_i_3 
       (.I0(\out[1544]_i_6_n_0 ),
        .I1(padder_out_1[548]),
        .I2(out[484]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1544]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1435]),
        .O(\out[1544]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1544]_i_4 
       (.I0(\out[1544]_i_9_n_0 ),
        .I1(padder_out_1[485]),
        .I2(out[421]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1544]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1372]),
        .O(\out[1544]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1544]_i_5 
       (.I0(\f_permutation_l_/round_in [1544]),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[1544]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1544]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[924] ),
        .I1(padder_out_1[228]),
        .I2(out[164]),
        .I3(\f_permutation_l_/out_reg_n_0_[284] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[604] ),
        .O(\out[1544]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1544]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[795] ),
        .I1(padder_out_1[99]),
        .I2(out[35]),
        .I3(\f_permutation_l_/out_reg_n_0_[155] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[475] ),
        .O(\out[1544]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1544]_i_8 
       (.I0(padder_out_1[419]),
        .I1(out[355]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1435]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1544]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[861] ),
        .I1(padder_out_1[165]),
        .I2(out[101]),
        .I3(\f_permutation_l_/out_reg_n_0_[221] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[541] ),
        .O(\out[1544]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1545]_i_1 
       (.I0(\f_permutation_l_/round_in [1181]),
        .I1(\out[1545]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[798] ),
        .I3(\out[1545]_i_4_n_0 ),
        .I4(\out[1545]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1545]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1545]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[733] ),
        .I1(padder_out_1[37]),
        .I2(\f_permutation_l_/out_reg_n_0_[1053] ),
        .I3(\f_permutation_l_/out_reg_n_0_[93] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[413] ),
        .O(\out[1545]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_11 
       (.I0(padder_out_1[357]),
        .I1(out[293]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1373]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_12 
       (.I0(padder_out_1[561]),
        .I1(out[497]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1545]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_13 
       (.I0(padder_out_1[305]),
        .I1(out[241]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1289]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1545]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[649] ),
        .I1(\f_permutation_l_/out_reg_n_0_[969] ),
        .I2(\f_permutation_l_/out_reg_n_0_[9] ),
        .I3(\f_permutation_l_/out_reg_n_0_[329] ),
        .O(\out[1545]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_15 
       (.I0(padder_out_1[496]),
        .I1(out[432]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1480]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1545]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[840] ),
        .I1(padder_out_1[176]),
        .I2(out[112]),
        .I3(\f_permutation_l_/out_reg_n_0_[200] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[520] ),
        .O(\out[1545]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_2 
       (.I0(padder_out_1[165]),
        .I1(out[101]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1181]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1545]_i_3 
       (.I0(\out[1545]_i_6_n_0 ),
        .I1(padder_out_1[549]),
        .I2(out[485]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1545]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1436]),
        .O(\out[1545]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1545]_i_4 
       (.I0(\out[1545]_i_9_n_0 ),
        .I1(padder_out_1[486]),
        .I2(out[422]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1545]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1373]),
        .O(\out[1545]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1545]_i_5 
       (.I0(\f_permutation_l_/round_in [1545]),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[1545]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1545]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[925] ),
        .I1(padder_out_1[229]),
        .I2(out[165]),
        .I3(\f_permutation_l_/out_reg_n_0_[285] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[605] ),
        .O(\out[1545]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1545]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[796] ),
        .I1(padder_out_1[100]),
        .I2(out[36]),
        .I3(\f_permutation_l_/out_reg_n_0_[156] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[476] ),
        .O(\out[1545]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1545]_i_8 
       (.I0(padder_out_1[420]),
        .I1(out[356]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1436]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1545]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[862] ),
        .I1(padder_out_1[166]),
        .I2(out[102]),
        .I3(\f_permutation_l_/out_reg_n_0_[222] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[542] ),
        .O(\out[1545]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1546]_i_1 
       (.I0(\f_permutation_l_/round_in [1182]),
        .I1(\out[1546]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[799] ),
        .I3(\out[1546]_i_4_n_0 ),
        .I4(\out[1546]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1546]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1546]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[734] ),
        .I1(padder_out_1[38]),
        .I2(\f_permutation_l_/out_reg_n_0_[1054] ),
        .I3(\f_permutation_l_/out_reg_n_0_[94] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[414] ),
        .O(\out[1546]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_11 
       (.I0(padder_out_1[358]),
        .I1(out[294]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1374]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_12 
       (.I0(padder_out_1[562]),
        .I1(out[498]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1546]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_13 
       (.I0(padder_out_1[306]),
        .I1(out[242]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1290]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1546]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[650] ),
        .I1(\f_permutation_l_/out_reg_n_0_[970] ),
        .I2(\f_permutation_l_/out_reg_n_0_[10] ),
        .I3(\f_permutation_l_/out_reg_n_0_[330] ),
        .O(\out[1546]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_15 
       (.I0(padder_out_1[497]),
        .I1(out[433]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1481]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1546]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[841] ),
        .I1(padder_out_1[177]),
        .I2(out[113]),
        .I3(\f_permutation_l_/out_reg_n_0_[201] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[521] ),
        .O(\out[1546]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_2 
       (.I0(padder_out_1[166]),
        .I1(out[102]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1182]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1546]_i_3 
       (.I0(\out[1546]_i_6_n_0 ),
        .I1(padder_out_1[550]),
        .I2(out[486]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1546]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1437]),
        .O(\out[1546]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1546]_i_4 
       (.I0(\out[1546]_i_9_n_0 ),
        .I1(padder_out_1[487]),
        .I2(out[423]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1546]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1374]),
        .O(\out[1546]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1546]_i_5 
       (.I0(\f_permutation_l_/round_in [1546]),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[1546]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1546]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[926] ),
        .I1(padder_out_1[230]),
        .I2(out[166]),
        .I3(\f_permutation_l_/out_reg_n_0_[286] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[606] ),
        .O(\out[1546]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1546]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[797] ),
        .I1(padder_out_1[101]),
        .I2(out[37]),
        .I3(\f_permutation_l_/out_reg_n_0_[157] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[477] ),
        .O(\out[1546]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1546]_i_8 
       (.I0(padder_out_1[421]),
        .I1(out[357]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1437]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1546]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[863] ),
        .I1(padder_out_1[167]),
        .I2(out[103]),
        .I3(\f_permutation_l_/out_reg_n_0_[223] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[543] ),
        .O(\out[1546]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1547]_i_1 
       (.I0(\f_permutation_l_/round_in [1183]),
        .I1(\out[1547]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[800] ),
        .I3(\out[1547]_i_4_n_0 ),
        .I4(\out[1547]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1547]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1547]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[735] ),
        .I1(padder_out_1[39]),
        .I2(\f_permutation_l_/out_reg_n_0_[1055] ),
        .I3(\f_permutation_l_/out_reg_n_0_[95] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[415] ),
        .O(\out[1547]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_11 
       (.I0(padder_out_1[359]),
        .I1(out[295]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1375]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_12 
       (.I0(padder_out_1[563]),
        .I1(out[499]),
        .I2(\out[1542]_i_8_n_0 ),
        .O(\f_permutation_l_/round_in [1547]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_13 
       (.I0(padder_out_1[307]),
        .I1(out[243]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1291]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1547]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[651] ),
        .I1(\f_permutation_l_/out_reg_n_0_[971] ),
        .I2(\f_permutation_l_/out_reg_n_0_[11] ),
        .I3(\f_permutation_l_/out_reg_n_0_[331] ),
        .O(\out[1547]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_15 
       (.I0(padder_out_1[498]),
        .I1(out[434]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1482]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1547]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[842] ),
        .I1(padder_out_1[178]),
        .I2(out[114]),
        .I3(\f_permutation_l_/out_reg_n_0_[202] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[522] ),
        .O(\out[1547]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_2 
       (.I0(padder_out_1[167]),
        .I1(out[103]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1183]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1547]_i_3 
       (.I0(\out[1547]_i_6_n_0 ),
        .I1(padder_out_1[551]),
        .I2(out[487]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1547]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1438]),
        .O(\out[1547]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1547]_i_4 
       (.I0(\out[1547]_i_9_n_0 ),
        .I1(padder_out_1[472]),
        .I2(out[408]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1547]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1375]),
        .O(\out[1547]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1547]_i_5 
       (.I0(\f_permutation_l_/round_in [1547]),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[1547]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1547]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[927] ),
        .I1(padder_out_1[231]),
        .I2(out[167]),
        .I3(\f_permutation_l_/out_reg_n_0_[287] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[607] ),
        .O(\out[1547]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1547]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[798] ),
        .I1(padder_out_1[102]),
        .I2(out[38]),
        .I3(\f_permutation_l_/out_reg_n_0_[158] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[478] ),
        .O(\out[1547]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1547]_i_8 
       (.I0(padder_out_1[422]),
        .I1(out[358]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1438]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1547]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[864] ),
        .I1(padder_out_1[152]),
        .I2(out[88]),
        .I3(\f_permutation_l_/out_reg_n_0_[224] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[544] ),
        .O(\out[1547]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1548]_i_1 
       (.I0(\f_permutation_l_/round_in [1184]),
        .I1(\out[1548]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[801] ),
        .I3(\out[1548]_i_4_n_0 ),
        .I4(\out[1548]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1548]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1548]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[736] ),
        .I1(padder_out_1[24]),
        .I2(\f_permutation_l_/out_reg_n_0_[1056] ),
        .I3(\f_permutation_l_/out_reg_n_0_[96] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[416] ),
        .O(\out[1548]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_11 
       (.I0(padder_out_1[344]),
        .I1(out[280]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1376]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_12 
       (.I0(padder_out_1[564]),
        .I1(out[500]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1548]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_13 
       (.I0(padder_out_1[308]),
        .I1(out[244]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1292]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1548]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[652] ),
        .I1(\f_permutation_l_/out_reg_n_0_[972] ),
        .I2(\f_permutation_l_/out_reg_n_0_[12] ),
        .I3(\f_permutation_l_/out_reg_n_0_[332] ),
        .O(\out[1548]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_15 
       (.I0(padder_out_1[499]),
        .I1(out[435]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1483]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1548]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[843] ),
        .I1(padder_out_1[179]),
        .I2(out[115]),
        .I3(\f_permutation_l_/out_reg_n_0_[203] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[523] ),
        .O(\out[1548]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_2 
       (.I0(padder_out_1[152]),
        .I1(out[88]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1184]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1548]_i_3 
       (.I0(\out[1548]_i_6_n_0 ),
        .I1(padder_out_1[536]),
        .I2(out[472]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1548]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1439]),
        .O(\out[1548]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1548]_i_4 
       (.I0(\out[1548]_i_9_n_0 ),
        .I1(padder_out_1[473]),
        .I2(out[409]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1548]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1376]),
        .O(\out[1548]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1548]_i_5 
       (.I0(\f_permutation_l_/round_in [1548]),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[1548]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1548]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[928] ),
        .I1(padder_out_1[216]),
        .I2(out[152]),
        .I3(\f_permutation_l_/out_reg_n_0_[288] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[608] ),
        .O(\out[1548]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1548]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[799] ),
        .I1(padder_out_1[103]),
        .I2(out[39]),
        .I3(\f_permutation_l_/out_reg_n_0_[159] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[479] ),
        .O(\out[1548]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1548]_i_8 
       (.I0(padder_out_1[423]),
        .I1(out[359]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1439]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1548]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[865] ),
        .I1(padder_out_1[153]),
        .I2(out[89]),
        .I3(\f_permutation_l_/out_reg_n_0_[225] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[545] ),
        .O(\out[1548]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1549]_i_1 
       (.I0(\f_permutation_l_/round_in [1185]),
        .I1(\out[1549]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[802] ),
        .I3(\out[1549]_i_4_n_0 ),
        .I4(\out[1549]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1549]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1549]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[737] ),
        .I1(padder_out_1[25]),
        .I2(\f_permutation_l_/out_reg_n_0_[1057] ),
        .I3(\f_permutation_l_/out_reg_n_0_[97] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[417] ),
        .O(\out[1549]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_11 
       (.I0(padder_out_1[345]),
        .I1(out[281]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1377]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_12 
       (.I0(padder_out_1[565]),
        .I1(out[501]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1549]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_13 
       (.I0(padder_out_1[309]),
        .I1(out[245]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1293]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1549]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[653] ),
        .I1(\f_permutation_l_/out_reg_n_0_[973] ),
        .I2(\f_permutation_l_/out_reg_n_0_[13] ),
        .I3(\f_permutation_l_/out_reg_n_0_[333] ),
        .O(\out[1549]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_15 
       (.I0(padder_out_1[500]),
        .I1(out[436]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1484]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1549]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[844] ),
        .I1(padder_out_1[180]),
        .I2(out[116]),
        .I3(\f_permutation_l_/out_reg_n_0_[204] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[524] ),
        .O(\out[1549]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_2 
       (.I0(padder_out_1[153]),
        .I1(out[89]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1185]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1549]_i_3 
       (.I0(\out[1549]_i_6_n_0 ),
        .I1(padder_out_1[537]),
        .I2(out[473]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1549]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1440]),
        .O(\out[1549]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1549]_i_4 
       (.I0(\out[1549]_i_9_n_0 ),
        .I1(padder_out_1[474]),
        .I2(out[410]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1549]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1377]),
        .O(\out[1549]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1549]_i_5 
       (.I0(\f_permutation_l_/round_in [1549]),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[1549]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1549]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[929] ),
        .I1(padder_out_1[217]),
        .I2(out[153]),
        .I3(\f_permutation_l_/out_reg_n_0_[289] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[609] ),
        .O(\out[1549]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1549]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[800] ),
        .I1(padder_out_1[88]),
        .I2(out[24]),
        .I3(\f_permutation_l_/out_reg_n_0_[160] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[480] ),
        .O(\out[1549]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1549]_i_8 
       (.I0(padder_out_1[408]),
        .I1(out[344]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1440]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1549]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[866] ),
        .I1(padder_out_1[154]),
        .I2(out[90]),
        .I3(\f_permutation_l_/out_reg_n_0_[226] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[546] ),
        .O(\out[1549]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[154]_i_1 
       (.I0(\out[1409]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[691] ),
        .I2(\out[154]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[216] ),
        .I4(\out[1540]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [154]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[154]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[625] ),
        .I1(\f_permutation_l_/round_in [1520]),
        .I2(\out[1563]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[154]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1550]_i_1 
       (.I0(\f_permutation_l_/round_in [1186]),
        .I1(\out[1550]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[803] ),
        .I3(\out[1550]_i_4_n_0 ),
        .I4(\out[1550]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1550]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1550]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[738] ),
        .I1(padder_out_1[26]),
        .I2(\f_permutation_l_/out_reg_n_0_[1058] ),
        .I3(\f_permutation_l_/out_reg_n_0_[98] ),
        .I4(\out[911]_i_4_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[418] ),
        .O(\out[1550]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_11 
       (.I0(padder_out_1[346]),
        .I1(out[282]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1378]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_12 
       (.I0(padder_out_1[566]),
        .I1(out[502]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1550]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_13 
       (.I0(padder_out_1[310]),
        .I1(out[246]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1294]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1550]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[654] ),
        .I1(\f_permutation_l_/out_reg_n_0_[974] ),
        .I2(\f_permutation_l_/out_reg_n_0_[14] ),
        .I3(\f_permutation_l_/out_reg_n_0_[334] ),
        .O(\out[1550]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_15 
       (.I0(padder_out_1[501]),
        .I1(out[437]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1485]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1550]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[845] ),
        .I1(padder_out_1[181]),
        .I2(out[117]),
        .I3(\f_permutation_l_/out_reg_n_0_[205] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[525] ),
        .O(\out[1550]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_2 
       (.I0(padder_out_1[154]),
        .I1(out[90]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1186]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1550]_i_3 
       (.I0(\out[1550]_i_6_n_0 ),
        .I1(padder_out_1[538]),
        .I2(out[474]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1550]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1441]),
        .O(\out[1550]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1550]_i_4 
       (.I0(\out[1550]_i_9_n_0 ),
        .I1(padder_out_1[475]),
        .I2(out[411]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1550]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1378]),
        .O(\out[1550]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1550]_i_5 
       (.I0(\f_permutation_l_/round_in [1550]),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[1550]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1550]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[930] ),
        .I1(padder_out_1[218]),
        .I2(out[154]),
        .I3(\f_permutation_l_/out_reg_n_0_[290] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[610] ),
        .O(\out[1550]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1550]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[801] ),
        .I1(padder_out_1[89]),
        .I2(out[25]),
        .I3(\f_permutation_l_/out_reg_n_0_[161] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[481] ),
        .O(\out[1550]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1550]_i_8 
       (.I0(padder_out_1[409]),
        .I1(out[345]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1441]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1550]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[867] ),
        .I1(padder_out_1[155]),
        .I2(out[91]),
        .I3(\f_permutation_l_/out_reg_n_0_[227] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[547] ),
        .O(\out[1550]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41BEBE41)) 
    \out[1551]_i_1 
       (.I0(\out[1551]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[804] ),
        .I2(\out[1551]_i_3_n_0 ),
        .I3(\out[1551]_i_4_n_0 ),
        .I4(\f_permutation_l_/rc [15]),
        .O(\f_permutation_l_/round_out [1551]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1551]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[868] ),
        .I1(padder_out_1[156]),
        .I2(out[92]),
        .I3(\f_permutation_l_/out_reg_n_0_[228] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[548] ),
        .O(\out[1551]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1551]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[739] ),
        .I1(padder_out_1[27]),
        .I2(\f_permutation_l_/out_reg_n_0_[1059] ),
        .I3(\f_permutation_l_/out_reg_n_0_[99] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[419] ),
        .O(\out[1551]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_12 
       (.I0(padder_out_1[347]),
        .I1(out[283]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1379]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_13 
       (.I0(padder_out_1[567]),
        .I1(out[503]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1551]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_14 
       (.I0(padder_out_1[311]),
        .I1(out[247]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1295]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1551]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[655] ),
        .I1(\f_permutation_l_/out_reg_n_0_[975] ),
        .I2(\f_permutation_l_/out_reg_n_0_[15] ),
        .I3(\f_permutation_l_/out_reg_n_0_[335] ),
        .O(\out[1551]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_16 
       (.I0(padder_out_1[502]),
        .I1(out[438]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1486]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1551]_i_17 
       (.I0(\f_permutation_l_/out_reg_n_0_[846] ),
        .I1(padder_out_1[182]),
        .I2(out[118]),
        .I3(\f_permutation_l_/out_reg_n_0_[206] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[526] ),
        .O(\out[1551]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \out[1551]_i_18 
       (.I0(\f_permutation_l_/i_reg_n_0_[15] ),
        .I1(\f_permutation_l_/i_reg_n_0_[14] ),
        .I2(\f_permutation_l_/i_reg_n_0_[2] ),
        .I3(\f_permutation_l_/p_0_in ),
        .O(\out[1551]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1551]_i_2 
       (.I0(\f_permutation_l_/round_in [1187]),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1571]),
        .I4(\out[1551]_i_9_n_0 ),
        .O(\out[1551]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1551]_i_3 
       (.I0(\out[1551]_i_10_n_0 ),
        .I1(padder_out_1[476]),
        .I2(out[412]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1551]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1379]),
        .O(\out[1551]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1551]_i_4 
       (.I0(\f_permutation_l_/round_in [1551]),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[1551]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1551]_i_5 
       (.I0(\f_permutation_l_/i_reg_n_0_ ),
        .I1(\out[1536]_i_6_n_0 ),
        .I2(\f_permutation_l_/i_reg_n_0_[17] ),
        .I3(\f_permutation_l_/i_reg_n_0_[1] ),
        .I4(\out[1543]_i_21_n_0 ),
        .I5(\out[1551]_i_18_n_0 ),
        .O(\f_permutation_l_/rc [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_6 
       (.I0(padder_out_1[410]),
        .I1(out[346]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1442]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1551]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[802] ),
        .I1(padder_out_1[90]),
        .I2(out[26]),
        .I3(\f_permutation_l_/out_reg_n_0_[162] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[482] ),
        .O(\out[1551]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1551]_i_8 
       (.I0(padder_out_1[539]),
        .I1(out[475]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1571]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1551]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[931] ),
        .I1(padder_out_1[219]),
        .I2(out[155]),
        .I3(\f_permutation_l_/out_reg_n_0_[291] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[611] ),
        .O(\out[1551]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1552]_i_1 
       (.I0(\f_permutation_l_/round_in [1188]),
        .I1(\out[1552]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[805] ),
        .I3(\out[1552]_i_4_n_0 ),
        .I4(\out[1552]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1552]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1552]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[740] ),
        .I1(padder_out_1[28]),
        .I2(\f_permutation_l_/out_reg_n_0_[1060] ),
        .I3(\f_permutation_l_/out_reg_n_0_[100] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[420] ),
        .O(\out[1552]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_11 
       (.I0(padder_out_1[348]),
        .I1(out[284]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1380]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_12 
       (.I0(padder_out_1[552]),
        .I1(out[488]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1552]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_13 
       (.I0(padder_out_1[296]),
        .I1(out[232]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1296]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1552]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[656] ),
        .I1(\f_permutation_l_/out_reg_n_0_[976] ),
        .I2(\f_permutation_l_/out_reg_n_0_[16] ),
        .I3(\f_permutation_l_/out_reg_n_0_[336] ),
        .O(\out[1552]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_15 
       (.I0(padder_out_1[503]),
        .I1(out[439]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1487]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1552]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[847] ),
        .I1(padder_out_1[183]),
        .I2(out[119]),
        .I3(\f_permutation_l_/out_reg_n_0_[207] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[527] ),
        .O(\out[1552]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_2 
       (.I0(padder_out_1[156]),
        .I1(out[92]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1188]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1552]_i_3 
       (.I0(\out[1552]_i_6_n_0 ),
        .I1(padder_out_1[540]),
        .I2(out[476]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1552]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1443]),
        .O(\out[1552]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1552]_i_4 
       (.I0(\out[1552]_i_9_n_0 ),
        .I1(padder_out_1[477]),
        .I2(out[413]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1552]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1380]),
        .O(\out[1552]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1552]_i_5 
       (.I0(\f_permutation_l_/round_in [1552]),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[1552]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1552]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[932] ),
        .I1(padder_out_1[220]),
        .I2(out[156]),
        .I3(\f_permutation_l_/out_reg_n_0_[292] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[612] ),
        .O(\out[1552]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1552]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[803] ),
        .I1(padder_out_1[91]),
        .I2(out[27]),
        .I3(\f_permutation_l_/out_reg_n_0_[163] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[483] ),
        .O(\out[1552]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1552]_i_8 
       (.I0(padder_out_1[411]),
        .I1(out[347]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1443]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1552]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[869] ),
        .I1(padder_out_1[157]),
        .I2(out[93]),
        .I3(\f_permutation_l_/out_reg_n_0_[229] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[549] ),
        .O(\out[1552]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1553]_i_1 
       (.I0(\f_permutation_l_/round_in [1189]),
        .I1(\out[1553]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[806] ),
        .I3(\out[1553]_i_4_n_0 ),
        .I4(\out[1553]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1553]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1553]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[741] ),
        .I1(padder_out_1[29]),
        .I2(\f_permutation_l_/out_reg_n_0_[1061] ),
        .I3(\f_permutation_l_/out_reg_n_0_[101] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[421] ),
        .O(\out[1553]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_11 
       (.I0(padder_out_1[349]),
        .I1(out[285]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1381]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_12 
       (.I0(padder_out_1[553]),
        .I1(out[489]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1553]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_13 
       (.I0(padder_out_1[297]),
        .I1(out[233]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1297]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1553]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[657] ),
        .I1(\f_permutation_l_/out_reg_n_0_[977] ),
        .I2(\f_permutation_l_/out_reg_n_0_[17] ),
        .I3(\f_permutation_l_/out_reg_n_0_[337] ),
        .O(\out[1553]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_15 
       (.I0(padder_out_1[488]),
        .I1(out[424]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1488]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1553]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[848] ),
        .I1(padder_out_1[168]),
        .I2(out[104]),
        .I3(\f_permutation_l_/out_reg_n_0_[208] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[528] ),
        .O(\out[1553]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_2 
       (.I0(padder_out_1[157]),
        .I1(out[93]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1189]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1553]_i_3 
       (.I0(\out[1553]_i_6_n_0 ),
        .I1(padder_out_1[541]),
        .I2(out[477]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1553]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1444]),
        .O(\out[1553]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1553]_i_4 
       (.I0(\out[1553]_i_9_n_0 ),
        .I1(padder_out_1[478]),
        .I2(out[414]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1553]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1381]),
        .O(\out[1553]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1553]_i_5 
       (.I0(\f_permutation_l_/round_in [1553]),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[1553]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1553]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[933] ),
        .I1(padder_out_1[221]),
        .I2(out[157]),
        .I3(\f_permutation_l_/out_reg_n_0_[293] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[613] ),
        .O(\out[1553]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1553]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[804] ),
        .I1(padder_out_1[92]),
        .I2(out[28]),
        .I3(\f_permutation_l_/out_reg_n_0_[164] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[484] ),
        .O(\out[1553]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1553]_i_8 
       (.I0(padder_out_1[412]),
        .I1(out[348]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1444]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1553]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[870] ),
        .I1(padder_out_1[158]),
        .I2(out[94]),
        .I3(\f_permutation_l_/out_reg_n_0_[230] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[550] ),
        .O(\out[1553]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1554]_i_1 
       (.I0(\f_permutation_l_/round_in [1190]),
        .I1(\out[1554]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[807] ),
        .I3(\out[1554]_i_4_n_0 ),
        .I4(\out[1554]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1554]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1554]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[742] ),
        .I1(padder_out_1[30]),
        .I2(\f_permutation_l_/out_reg_n_0_[1062] ),
        .I3(\f_permutation_l_/out_reg_n_0_[102] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[422] ),
        .O(\out[1554]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_11 
       (.I0(padder_out_1[350]),
        .I1(out[286]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1382]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_12 
       (.I0(padder_out_1[554]),
        .I1(out[490]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1554]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_13 
       (.I0(padder_out_1[298]),
        .I1(out[234]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1298]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1554]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[658] ),
        .I1(\f_permutation_l_/out_reg_n_0_[978] ),
        .I2(\f_permutation_l_/out_reg_n_0_[18] ),
        .I3(\f_permutation_l_/out_reg_n_0_[338] ),
        .O(\out[1554]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_15 
       (.I0(padder_out_1[489]),
        .I1(out[425]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1489]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1554]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[849] ),
        .I1(padder_out_1[169]),
        .I2(out[105]),
        .I3(\f_permutation_l_/out_reg_n_0_[209] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[529] ),
        .O(\out[1554]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_2 
       (.I0(padder_out_1[158]),
        .I1(out[94]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1190]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1554]_i_3 
       (.I0(\out[1554]_i_6_n_0 ),
        .I1(padder_out_1[542]),
        .I2(out[478]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1554]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1445]),
        .O(\out[1554]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1554]_i_4 
       (.I0(\out[1554]_i_9_n_0 ),
        .I1(padder_out_1[479]),
        .I2(out[415]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1554]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1382]),
        .O(\out[1554]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1554]_i_5 
       (.I0(\f_permutation_l_/round_in [1554]),
        .I1(\f_permutation_l_/round_in [1298]),
        .I2(\out[1554]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[1554]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1554]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[934] ),
        .I1(padder_out_1[222]),
        .I2(out[158]),
        .I3(\f_permutation_l_/out_reg_n_0_[294] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[614] ),
        .O(\out[1554]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1554]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[805] ),
        .I1(padder_out_1[93]),
        .I2(out[29]),
        .I3(\f_permutation_l_/out_reg_n_0_[165] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[485] ),
        .O(\out[1554]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1554]_i_8 
       (.I0(padder_out_1[413]),
        .I1(out[349]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1445]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1554]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[871] ),
        .I1(padder_out_1[159]),
        .I2(out[95]),
        .I3(\f_permutation_l_/out_reg_n_0_[231] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[551] ),
        .O(\out[1554]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1555]_i_1 
       (.I0(\f_permutation_l_/round_in [1191]),
        .I1(\out[1555]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[808] ),
        .I3(\out[1555]_i_4_n_0 ),
        .I4(\out[1555]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1555]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1555]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[743] ),
        .I1(padder_out_1[31]),
        .I2(\f_permutation_l_/out_reg_n_0_[1063] ),
        .I3(\f_permutation_l_/out_reg_n_0_[103] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[423] ),
        .O(\out[1555]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_11 
       (.I0(padder_out_1[351]),
        .I1(out[287]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1383]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_12 
       (.I0(padder_out_1[555]),
        .I1(out[491]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1555]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_13 
       (.I0(padder_out_1[299]),
        .I1(out[235]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1299]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1555]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[659] ),
        .I1(\f_permutation_l_/out_reg_n_0_[979] ),
        .I2(\f_permutation_l_/out_reg_n_0_[19] ),
        .I3(\f_permutation_l_/out_reg_n_0_[339] ),
        .O(\out[1555]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_15 
       (.I0(padder_out_1[490]),
        .I1(out[426]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1490]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1555]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[850] ),
        .I1(padder_out_1[170]),
        .I2(out[106]),
        .I3(\f_permutation_l_/out_reg_n_0_[210] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[530] ),
        .O(\out[1555]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_2 
       (.I0(padder_out_1[159]),
        .I1(out[95]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1191]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1555]_i_3 
       (.I0(\out[1555]_i_6_n_0 ),
        .I1(padder_out_1[543]),
        .I2(out[479]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1555]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1446]),
        .O(\out[1555]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1555]_i_4 
       (.I0(\out[1555]_i_9_n_0 ),
        .I1(padder_out_1[464]),
        .I2(out[400]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1555]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1383]),
        .O(\out[1555]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1555]_i_5 
       (.I0(\f_permutation_l_/round_in [1555]),
        .I1(\f_permutation_l_/round_in [1299]),
        .I2(\out[1555]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[1555]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1555]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[935] ),
        .I1(padder_out_1[223]),
        .I2(out[159]),
        .I3(\f_permutation_l_/out_reg_n_0_[295] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[615] ),
        .O(\out[1555]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1555]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[806] ),
        .I1(padder_out_1[94]),
        .I2(out[30]),
        .I3(\f_permutation_l_/out_reg_n_0_[166] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[486] ),
        .O(\out[1555]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1555]_i_8 
       (.I0(padder_out_1[414]),
        .I1(out[350]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1446]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1555]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[872] ),
        .I1(padder_out_1[144]),
        .I2(out[80]),
        .I3(\f_permutation_l_/out_reg_n_0_[232] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[552] ),
        .O(\out[1555]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1556]_i_1 
       (.I0(\f_permutation_l_/round_in [1192]),
        .I1(\out[1556]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[809] ),
        .I3(\out[1556]_i_4_n_0 ),
        .I4(\out[1556]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1556]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1556]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[873] ),
        .I1(padder_out_1[145]),
        .I2(out[81]),
        .I3(\f_permutation_l_/out_reg_n_0_[233] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[553] ),
        .O(\out[1556]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1556]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[744] ),
        .I1(padder_out_1[16]),
        .I2(\f_permutation_l_/out_reg_n_0_[1064] ),
        .I3(\f_permutation_l_/out_reg_n_0_[104] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[424] ),
        .O(\out[1556]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1556]_i_12 
       (.I0(padder_out_1[336]),
        .I1(out[272]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1384]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1556]_i_13 
       (.I0(padder_out_1[300]),
        .I1(out[236]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1300]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1556]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[660] ),
        .I1(\f_permutation_l_/out_reg_n_0_[980] ),
        .I2(\f_permutation_l_/out_reg_n_0_[20] ),
        .I3(\f_permutation_l_/out_reg_n_0_[340] ),
        .O(\out[1556]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1556]_i_15 
       (.I0(padder_out_1[491]),
        .I1(out[427]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1491]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1556]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[851] ),
        .I1(padder_out_1[171]),
        .I2(out[107]),
        .I3(\f_permutation_l_/out_reg_n_0_[211] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[531] ),
        .O(\out[1556]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1556]_i_2 
       (.I0(padder_out_1[144]),
        .I1(out[80]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1192]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1556]_i_3 
       (.I0(\out[1556]_i_6_n_0 ),
        .I1(padder_out_1[528]),
        .I2(out[464]),
        .I3(\out[1556]_i_7_n_0 ),
        .I4(\out[1556]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1447]),
        .O(\out[1556]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1556]_i_4 
       (.I0(\out[1556]_i_10_n_0 ),
        .I1(padder_out_1[465]),
        .I2(out[401]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1556]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1384]),
        .O(\out[1556]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1556]_i_5 
       (.I0(\f_permutation_l_/round_in [1556]),
        .I1(\f_permutation_l_/round_in [1300]),
        .I2(\out[1556]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[1556]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1556]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[936] ),
        .I1(padder_out_1[208]),
        .I2(out[144]),
        .I3(\f_permutation_l_/out_reg_n_0_[296] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[616] ),
        .O(\out[1556]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1556]_i_7 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1556]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1556]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[807] ),
        .I1(padder_out_1[95]),
        .I2(out[31]),
        .I3(\f_permutation_l_/out_reg_n_0_[167] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[487] ),
        .O(\out[1556]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1556]_i_9 
       (.I0(padder_out_1[415]),
        .I1(out[351]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1447]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1557]_i_1 
       (.I0(\f_permutation_l_/round_in [1193]),
        .I1(\out[1557]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[810] ),
        .I3(\out[1557]_i_4_n_0 ),
        .I4(\out[1557]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1557]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1557]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[745] ),
        .I1(padder_out_1[17]),
        .I2(\f_permutation_l_/out_reg_n_0_[1065] ),
        .I3(\f_permutation_l_/out_reg_n_0_[105] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[425] ),
        .O(\out[1557]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1557]_i_11 
       (.I0(padder_out_1[337]),
        .I1(out[273]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1385]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1557]_i_12 
       (.I0(padder_out_1[301]),
        .I1(out[237]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1301]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1557]_i_13 
       (.I0(\f_permutation_l_/out_reg_n_0_[661] ),
        .I1(\f_permutation_l_/out_reg_n_0_[981] ),
        .I2(\f_permutation_l_/out_reg_n_0_[21] ),
        .I3(\f_permutation_l_/out_reg_n_0_[341] ),
        .O(\out[1557]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1557]_i_14 
       (.I0(padder_out_1[492]),
        .I1(out[428]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1492]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1557]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[852] ),
        .I1(padder_out_1[172]),
        .I2(out[108]),
        .I3(\f_permutation_l_/out_reg_n_0_[212] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[532] ),
        .O(\out[1557]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1557]_i_2 
       (.I0(padder_out_1[145]),
        .I1(out[81]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1193]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1557]_i_3 
       (.I0(\out[1557]_i_6_n_0 ),
        .I1(padder_out_1[529]),
        .I2(out[465]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1557]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1448]),
        .O(\out[1557]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1557]_i_4 
       (.I0(\out[1557]_i_9_n_0 ),
        .I1(padder_out_1[466]),
        .I2(out[402]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1557]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1385]),
        .O(\out[1557]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1557]_i_5 
       (.I0(\f_permutation_l_/round_in [1557]),
        .I1(\f_permutation_l_/round_in [1301]),
        .I2(\out[1557]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[1557]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1557]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[937] ),
        .I1(padder_out_1[209]),
        .I2(out[145]),
        .I3(\f_permutation_l_/out_reg_n_0_[297] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[617] ),
        .O(\out[1557]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1557]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[808] ),
        .I1(padder_out_1[80]),
        .I2(out[16]),
        .I3(\f_permutation_l_/out_reg_n_0_[168] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[488] ),
        .O(\out[1557]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1557]_i_8 
       (.I0(padder_out_1[400]),
        .I1(out[336]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1448]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1557]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[874] ),
        .I1(padder_out_1[146]),
        .I2(out[82]),
        .I3(\f_permutation_l_/out_reg_n_0_[234] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[554] ),
        .O(\out[1557]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1558]_i_1 
       (.I0(\f_permutation_l_/round_in [1194]),
        .I1(\out[1558]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[811] ),
        .I3(\out[1558]_i_4_n_0 ),
        .I4(\out[1558]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1558]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1558]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[746] ),
        .I1(padder_out_1[18]),
        .I2(\f_permutation_l_/out_reg_n_0_[1066] ),
        .I3(\f_permutation_l_/out_reg_n_0_[106] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[426] ),
        .O(\out[1558]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1558]_i_11 
       (.I0(padder_out_1[338]),
        .I1(out[274]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1386]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1558]_i_12 
       (.I0(padder_out_1[558]),
        .I1(out[494]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1558]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1558]_i_13 
       (.I0(padder_out_1[302]),
        .I1(out[238]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1302]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1558]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[662] ),
        .I1(\f_permutation_l_/out_reg_n_0_[982] ),
        .I2(\f_permutation_l_/out_reg_n_0_[22] ),
        .I3(\f_permutation_l_/out_reg_n_0_[342] ),
        .O(\out[1558]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1558]_i_2 
       (.I0(padder_out_1[146]),
        .I1(out[82]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1194]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1558]_i_3 
       (.I0(\out[1558]_i_6_n_0 ),
        .I1(padder_out_1[530]),
        .I2(out[466]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1558]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1449]),
        .O(\out[1558]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1558]_i_4 
       (.I0(\out[1558]_i_9_n_0 ),
        .I1(padder_out_1[467]),
        .I2(out[403]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1558]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1386]),
        .O(\out[1558]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1558]_i_5 
       (.I0(\f_permutation_l_/round_in [1558]),
        .I1(\out[1536]_i_14_n_0 ),
        .I2(\f_permutation_l_/round_in [1493]),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[1558]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1558]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[938] ),
        .I1(padder_out_1[210]),
        .I2(out[146]),
        .I3(\f_permutation_l_/out_reg_n_0_[298] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[618] ),
        .O(\out[1558]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1558]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[809] ),
        .I1(padder_out_1[81]),
        .I2(out[17]),
        .I3(\f_permutation_l_/out_reg_n_0_[169] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[489] ),
        .O(\out[1558]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1558]_i_8 
       (.I0(padder_out_1[401]),
        .I1(out[337]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1449]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1558]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[875] ),
        .I1(padder_out_1[147]),
        .I2(out[83]),
        .I3(\f_permutation_l_/out_reg_n_0_[235] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[555] ),
        .O(\out[1558]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1559]_i_1 
       (.I0(\f_permutation_l_/round_in [1195]),
        .I1(\out[1559]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[812] ),
        .I3(\out[1559]_i_4_n_0 ),
        .I4(\out[1559]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1559]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1559]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[747] ),
        .I1(padder_out_1[19]),
        .I2(\f_permutation_l_/out_reg_n_0_[1067] ),
        .I3(\f_permutation_l_/out_reg_n_0_[107] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[427] ),
        .O(\out[1559]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_11 
       (.I0(padder_out_1[339]),
        .I1(out[275]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1387]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_12 
       (.I0(padder_out_1[559]),
        .I1(out[495]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1559]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_13 
       (.I0(padder_out_1[494]),
        .I1(out[430]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1494]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_14 
       (.I0(padder_out_1[303]),
        .I1(out[239]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1303]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1559]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[663] ),
        .I1(\f_permutation_l_/out_reg_n_0_[983] ),
        .I2(\f_permutation_l_/out_reg_n_0_[23] ),
        .I3(\f_permutation_l_/out_reg_n_0_[343] ),
        .O(\out[1559]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_2 
       (.I0(padder_out_1[147]),
        .I1(out[83]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1195]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1559]_i_3 
       (.I0(\out[1559]_i_6_n_0 ),
        .I1(padder_out_1[531]),
        .I2(out[467]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1559]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1450]),
        .O(\out[1559]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1559]_i_4 
       (.I0(\out[1559]_i_9_n_0 ),
        .I1(padder_out_1[468]),
        .I2(out[404]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1559]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1387]),
        .O(\out[1559]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1559]_i_5 
       (.I0(\f_permutation_l_/round_in [1559]),
        .I1(\f_permutation_l_/round_in [1494]),
        .I2(\out[1537]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[1559]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1559]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[939] ),
        .I1(padder_out_1[211]),
        .I2(out[147]),
        .I3(\f_permutation_l_/out_reg_n_0_[299] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[619] ),
        .O(\out[1559]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1559]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[810] ),
        .I1(padder_out_1[82]),
        .I2(out[18]),
        .I3(\f_permutation_l_/out_reg_n_0_[170] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[490] ),
        .O(\out[1559]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1559]_i_8 
       (.I0(padder_out_1[402]),
        .I1(out[338]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1450]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1559]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[876] ),
        .I1(padder_out_1[148]),
        .I2(out[84]),
        .I3(\f_permutation_l_/out_reg_n_0_[236] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[556] ),
        .O(\out[1559]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[155]_i_1 
       (.I0(\out[1410]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[692] ),
        .I2(\out[155]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[217] ),
        .I4(\out[1541]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [155]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[155]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[626] ),
        .I1(\f_permutation_l_/round_in [1521]),
        .I2(\out[1564]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[155]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1560]_i_1 
       (.I0(\f_permutation_l_/round_in [1196]),
        .I1(\out[1560]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[813] ),
        .I3(\out[1560]_i_4_n_0 ),
        .I4(\out[1560]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1560]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1560]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[748] ),
        .I1(padder_out_1[20]),
        .I2(\f_permutation_l_/out_reg_n_0_[1068] ),
        .I3(\f_permutation_l_/out_reg_n_0_[108] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[428] ),
        .O(\out[1560]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_11 
       (.I0(padder_out_1[340]),
        .I1(out[276]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1388]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_12 
       (.I0(padder_out_1[544]),
        .I1(out[480]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1560]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_13 
       (.I0(padder_out_1[495]),
        .I1(out[431]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1495]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_14 
       (.I0(padder_out_1[288]),
        .I1(out[224]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1304]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1560]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[664] ),
        .I1(\f_permutation_l_/out_reg_n_0_[984] ),
        .I2(\f_permutation_l_/out_reg_n_0_[24] ),
        .I3(\f_permutation_l_/out_reg_n_0_[344] ),
        .O(\out[1560]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_2 
       (.I0(padder_out_1[148]),
        .I1(out[84]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1196]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1560]_i_3 
       (.I0(\out[1560]_i_6_n_0 ),
        .I1(padder_out_1[532]),
        .I2(out[468]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1560]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1451]),
        .O(\out[1560]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1560]_i_4 
       (.I0(\out[1560]_i_9_n_0 ),
        .I1(padder_out_1[469]),
        .I2(out[405]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1560]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1388]),
        .O(\out[1560]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1560]_i_5 
       (.I0(\f_permutation_l_/round_in [1560]),
        .I1(\f_permutation_l_/round_in [1495]),
        .I2(\out[1538]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[1560]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1560]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[940] ),
        .I1(padder_out_1[212]),
        .I2(out[148]),
        .I3(\f_permutation_l_/out_reg_n_0_[300] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[620] ),
        .O(\out[1560]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1560]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[811] ),
        .I1(padder_out_1[83]),
        .I2(out[19]),
        .I3(\f_permutation_l_/out_reg_n_0_[171] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[491] ),
        .O(\out[1560]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1560]_i_8 
       (.I0(padder_out_1[403]),
        .I1(out[339]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1451]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1560]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[877] ),
        .I1(padder_out_1[149]),
        .I2(out[85]),
        .I3(\f_permutation_l_/out_reg_n_0_[237] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[557] ),
        .O(\out[1560]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1561]_i_1 
       (.I0(\f_permutation_l_/round_in [1197]),
        .I1(\out[1561]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[814] ),
        .I3(\out[1561]_i_4_n_0 ),
        .I4(\out[1561]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1561]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1561]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[749] ),
        .I1(padder_out_1[21]),
        .I2(\f_permutation_l_/out_reg_n_0_[1069] ),
        .I3(\f_permutation_l_/out_reg_n_0_[109] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[429] ),
        .O(\out[1561]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1561]_i_11 
       (.I0(padder_out_1[341]),
        .I1(out[277]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1389]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1561]_i_12 
       (.I0(padder_out_1[545]),
        .I1(out[481]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1561]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1561]_i_13 
       (.I0(padder_out_1[289]),
        .I1(out[225]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1305]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1561]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[665] ),
        .I1(\f_permutation_l_/out_reg_n_0_[985] ),
        .I2(\f_permutation_l_/out_reg_n_0_[25] ),
        .I3(\f_permutation_l_/out_reg_n_0_[345] ),
        .O(\out[1561]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1561]_i_2 
       (.I0(padder_out_1[149]),
        .I1(out[85]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1197]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1561]_i_3 
       (.I0(\out[1561]_i_6_n_0 ),
        .I1(padder_out_1[533]),
        .I2(out[469]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1561]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1452]),
        .O(\out[1561]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1561]_i_4 
       (.I0(\out[1561]_i_9_n_0 ),
        .I1(padder_out_1[470]),
        .I2(out[406]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1561]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1389]),
        .O(\out[1561]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1561]_i_5 
       (.I0(\f_permutation_l_/round_in [1561]),
        .I1(\f_permutation_l_/round_in [1496]),
        .I2(\out[1539]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[1561]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1561]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[941] ),
        .I1(padder_out_1[213]),
        .I2(out[149]),
        .I3(\f_permutation_l_/out_reg_n_0_[301] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[621] ),
        .O(\out[1561]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1561]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[812] ),
        .I1(padder_out_1[84]),
        .I2(out[20]),
        .I3(\f_permutation_l_/out_reg_n_0_[172] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[492] ),
        .O(\out[1561]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1561]_i_8 
       (.I0(padder_out_1[404]),
        .I1(out[340]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1452]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1561]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[878] ),
        .I1(padder_out_1[150]),
        .I2(out[86]),
        .I3(\f_permutation_l_/out_reg_n_0_[238] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[558] ),
        .O(\out[1561]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1562]_i_1 
       (.I0(\f_permutation_l_/round_in [1198]),
        .I1(\out[1562]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[815] ),
        .I3(\out[1562]_i_4_n_0 ),
        .I4(\out[1562]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1562]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1562]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[750] ),
        .I1(padder_out_1[22]),
        .I2(\f_permutation_l_/out_reg_n_0_[1070] ),
        .I3(\f_permutation_l_/out_reg_n_0_[110] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[430] ),
        .O(\out[1562]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_11 
       (.I0(padder_out_1[342]),
        .I1(out[278]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1390]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_12 
       (.I0(padder_out_1[546]),
        .I1(out[482]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1562]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_13 
       (.I0(padder_out_1[481]),
        .I1(out[417]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1497]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_14 
       (.I0(padder_out_1[290]),
        .I1(out[226]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1306]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1562]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[666] ),
        .I1(\f_permutation_l_/out_reg_n_0_[986] ),
        .I2(\f_permutation_l_/out_reg_n_0_[26] ),
        .I3(\f_permutation_l_/out_reg_n_0_[346] ),
        .O(\out[1562]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_2 
       (.I0(padder_out_1[150]),
        .I1(out[86]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1198]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1562]_i_3 
       (.I0(\out[1562]_i_6_n_0 ),
        .I1(padder_out_1[534]),
        .I2(out[470]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1562]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1453]),
        .O(\out[1562]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1562]_i_4 
       (.I0(\out[1562]_i_9_n_0 ),
        .I1(padder_out_1[471]),
        .I2(out[407]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1562]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1390]),
        .O(\out[1562]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1562]_i_5 
       (.I0(\f_permutation_l_/round_in [1562]),
        .I1(\f_permutation_l_/round_in [1497]),
        .I2(\out[1540]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[1562]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1562]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[942] ),
        .I1(padder_out_1[214]),
        .I2(out[150]),
        .I3(\f_permutation_l_/out_reg_n_0_[302] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[622] ),
        .O(\out[1562]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1562]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[813] ),
        .I1(padder_out_1[85]),
        .I2(out[21]),
        .I3(\f_permutation_l_/out_reg_n_0_[173] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[493] ),
        .O(\out[1562]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1562]_i_8 
       (.I0(padder_out_1[405]),
        .I1(out[341]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1453]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1562]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[879] ),
        .I1(padder_out_1[151]),
        .I2(out[87]),
        .I3(\f_permutation_l_/out_reg_n_0_[239] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[559] ),
        .O(\out[1562]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1563]_i_1 
       (.I0(\f_permutation_l_/round_in [1199]),
        .I1(\out[1563]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[816] ),
        .I3(\out[1563]_i_4_n_0 ),
        .I4(\out[1563]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1563]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1563]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[751] ),
        .I1(padder_out_1[23]),
        .I2(\f_permutation_l_/out_reg_n_0_[1071] ),
        .I3(\f_permutation_l_/out_reg_n_0_[111] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[431] ),
        .O(\out[1563]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1563]_i_11 
       (.I0(padder_out_1[343]),
        .I1(out[279]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1391]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1563]_i_12 
       (.I0(padder_out_1[482]),
        .I1(out[418]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1498]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1563]_i_13 
       (.I0(padder_out_1[291]),
        .I1(out[227]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1307]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1563]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[667] ),
        .I1(\f_permutation_l_/out_reg_n_0_[987] ),
        .I2(\f_permutation_l_/out_reg_n_0_[27] ),
        .I3(\f_permutation_l_/out_reg_n_0_[347] ),
        .O(\out[1563]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1563]_i_2 
       (.I0(padder_out_1[151]),
        .I1(out[87]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1199]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1563]_i_3 
       (.I0(\out[1563]_i_6_n_0 ),
        .I1(padder_out_1[535]),
        .I2(out[471]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1563]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1454]),
        .O(\out[1563]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1563]_i_4 
       (.I0(\out[1563]_i_9_n_0 ),
        .I1(padder_out_1[456]),
        .I2(out[392]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1563]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1391]),
        .O(\out[1563]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1563]_i_5 
       (.I0(\f_permutation_l_/round_in [1563]),
        .I1(\f_permutation_l_/round_in [1498]),
        .I2(\out[1541]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[1563]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1563]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[943] ),
        .I1(padder_out_1[215]),
        .I2(out[151]),
        .I3(\f_permutation_l_/out_reg_n_0_[303] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[623] ),
        .O(\out[1563]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1563]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[814] ),
        .I1(padder_out_1[86]),
        .I2(out[22]),
        .I3(\f_permutation_l_/out_reg_n_0_[174] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[494] ),
        .O(\out[1563]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1563]_i_8 
       (.I0(padder_out_1[406]),
        .I1(out[342]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1454]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1563]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[880] ),
        .I1(padder_out_1[136]),
        .I2(out[72]),
        .I3(\f_permutation_l_/out_reg_n_0_[240] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[560] ),
        .O(\out[1563]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1564]_i_1 
       (.I0(\f_permutation_l_/round_in [1200]),
        .I1(\out[1564]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[817] ),
        .I3(\out[1564]_i_4_n_0 ),
        .I4(\out[1564]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1564]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1564]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[752] ),
        .I1(padder_out_1[8]),
        .I2(\f_permutation_l_/out_reg_n_0_[1072] ),
        .I3(\f_permutation_l_/out_reg_n_0_[112] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[432] ),
        .O(\out[1564]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_11 
       (.I0(padder_out_1[328]),
        .I1(out[264]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1392]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_12 
       (.I0(padder_out_1[548]),
        .I1(out[484]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1564]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_13 
       (.I0(padder_out_1[483]),
        .I1(out[419]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1499]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_14 
       (.I0(padder_out_1[292]),
        .I1(out[228]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1308]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1564]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[668] ),
        .I1(\f_permutation_l_/out_reg_n_0_[988] ),
        .I2(\f_permutation_l_/out_reg_n_0_[28] ),
        .I3(\f_permutation_l_/out_reg_n_0_[348] ),
        .O(\out[1564]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_2 
       (.I0(padder_out_1[136]),
        .I1(out[72]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1200]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1564]_i_3 
       (.I0(\out[1564]_i_6_n_0 ),
        .I1(padder_out_1[520]),
        .I2(out[456]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1564]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1455]),
        .O(\out[1564]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1564]_i_4 
       (.I0(\out[1564]_i_9_n_0 ),
        .I1(padder_out_1[457]),
        .I2(out[393]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1564]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1392]),
        .O(\out[1564]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1564]_i_5 
       (.I0(\f_permutation_l_/round_in [1564]),
        .I1(\f_permutation_l_/round_in [1499]),
        .I2(\out[1542]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[1564]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1564]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[944] ),
        .I1(padder_out_1[200]),
        .I2(out[136]),
        .I3(\f_permutation_l_/out_reg_n_0_[304] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[624] ),
        .O(\out[1564]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1564]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[815] ),
        .I1(padder_out_1[87]),
        .I2(out[23]),
        .I3(\f_permutation_l_/out_reg_n_0_[175] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[495] ),
        .O(\out[1564]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1564]_i_8 
       (.I0(padder_out_1[407]),
        .I1(out[343]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1455]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1564]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[881] ),
        .I1(padder_out_1[137]),
        .I2(out[73]),
        .I3(\f_permutation_l_/out_reg_n_0_[241] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[561] ),
        .O(\out[1564]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1565]_i_1 
       (.I0(\f_permutation_l_/round_in [1201]),
        .I1(\out[1565]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[818] ),
        .I3(\out[1565]_i_4_n_0 ),
        .I4(\out[1565]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1565]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1565]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[753] ),
        .I1(padder_out_1[9]),
        .I2(\f_permutation_l_/out_reg_n_0_[1073] ),
        .I3(\f_permutation_l_/out_reg_n_0_[113] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[433] ),
        .O(\out[1565]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_11 
       (.I0(padder_out_1[329]),
        .I1(out[265]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1393]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_12 
       (.I0(padder_out_1[549]),
        .I1(out[485]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1565]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_13 
       (.I0(padder_out_1[484]),
        .I1(out[420]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1500]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_14 
       (.I0(padder_out_1[293]),
        .I1(out[229]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1309]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1565]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[669] ),
        .I1(\f_permutation_l_/out_reg_n_0_[989] ),
        .I2(\f_permutation_l_/out_reg_n_0_[29] ),
        .I3(\f_permutation_l_/out_reg_n_0_[349] ),
        .O(\out[1565]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_2 
       (.I0(padder_out_1[137]),
        .I1(out[73]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1201]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1565]_i_3 
       (.I0(\out[1565]_i_6_n_0 ),
        .I1(padder_out_1[521]),
        .I2(out[457]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1565]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1456]),
        .O(\out[1565]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1565]_i_4 
       (.I0(\out[1565]_i_9_n_0 ),
        .I1(padder_out_1[458]),
        .I2(out[394]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1565]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1393]),
        .O(\out[1565]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1565]_i_5 
       (.I0(\f_permutation_l_/round_in [1565]),
        .I1(\f_permutation_l_/round_in [1500]),
        .I2(\out[1543]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[1565]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1565]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[945] ),
        .I1(padder_out_1[201]),
        .I2(out[137]),
        .I3(\f_permutation_l_/out_reg_n_0_[305] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[625] ),
        .O(\out[1565]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1565]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[816] ),
        .I1(padder_out_1[72]),
        .I2(out[8]),
        .I3(\f_permutation_l_/out_reg_n_0_[176] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[496] ),
        .O(\out[1565]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1565]_i_8 
       (.I0(padder_out_1[392]),
        .I1(out[328]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1456]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1565]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[882] ),
        .I1(padder_out_1[138]),
        .I2(out[74]),
        .I3(\f_permutation_l_/out_reg_n_0_[242] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[562] ),
        .O(\out[1565]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1566]_i_1 
       (.I0(\f_permutation_l_/round_in [1202]),
        .I1(\out[1566]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[819] ),
        .I3(\out[1566]_i_4_n_0 ),
        .I4(\out[1566]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1566]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1566]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[754] ),
        .I1(padder_out_1[10]),
        .I2(\f_permutation_l_/out_reg_n_0_[1074] ),
        .I3(\f_permutation_l_/out_reg_n_0_[114] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[434] ),
        .O(\out[1566]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1566]_i_11 
       (.I0(padder_out_1[330]),
        .I1(out[266]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1394]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1566]_i_12 
       (.I0(padder_out_1[550]),
        .I1(out[486]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1566]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1566]_i_13 
       (.I0(padder_out_1[294]),
        .I1(out[230]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1310]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1566]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[670] ),
        .I1(\f_permutation_l_/out_reg_n_0_[990] ),
        .I2(\f_permutation_l_/out_reg_n_0_[30] ),
        .I3(\f_permutation_l_/out_reg_n_0_[350] ),
        .O(\out[1566]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1566]_i_2 
       (.I0(padder_out_1[138]),
        .I1(out[74]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1202]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1566]_i_3 
       (.I0(\out[1566]_i_6_n_0 ),
        .I1(padder_out_1[522]),
        .I2(out[458]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1566]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1457]),
        .O(\out[1566]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1566]_i_4 
       (.I0(\out[1566]_i_9_n_0 ),
        .I1(padder_out_1[459]),
        .I2(out[395]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1566]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1394]),
        .O(\out[1566]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1566]_i_5 
       (.I0(\f_permutation_l_/round_in [1566]),
        .I1(\f_permutation_l_/round_in [1501]),
        .I2(\out[1544]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[1566]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1566]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[946] ),
        .I1(padder_out_1[202]),
        .I2(out[138]),
        .I3(\f_permutation_l_/out_reg_n_0_[306] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[626] ),
        .O(\out[1566]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1566]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[817] ),
        .I1(padder_out_1[73]),
        .I2(out[9]),
        .I3(\f_permutation_l_/out_reg_n_0_[177] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[497] ),
        .O(\out[1566]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1566]_i_8 
       (.I0(padder_out_1[393]),
        .I1(out[329]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1457]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1566]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[883] ),
        .I1(padder_out_1[139]),
        .I2(out[75]),
        .I3(\f_permutation_l_/out_reg_n_0_[243] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[563] ),
        .O(\out[1566]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41BEBE41)) 
    \out[1567]_i_1 
       (.I0(\out[1567]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[820] ),
        .I2(\out[1567]_i_3_n_0 ),
        .I3(\out[1567]_i_4_n_0 ),
        .I4(\f_permutation_l_/rc [31]),
        .O(\f_permutation_l_/round_out [1567]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1567]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[884] ),
        .I1(padder_out_1[140]),
        .I2(out[76]),
        .I3(\f_permutation_l_/out_reg_n_0_[244] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[564] ),
        .O(\out[1567]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1567]_i_11 
       (.I0(\f_permutation_l_/out_reg_n_0_[755] ),
        .I1(padder_out_1[11]),
        .I2(\f_permutation_l_/out_reg_n_0_[1075] ),
        .I3(\f_permutation_l_/out_reg_n_0_[115] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[435] ),
        .O(\out[1567]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_12 
       (.I0(padder_out_1[331]),
        .I1(out[267]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1395]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_13 
       (.I0(padder_out_1[551]),
        .I1(out[487]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1567]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_14 
       (.I0(padder_out_1[486]),
        .I1(out[422]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1502]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_15 
       (.I0(padder_out_1[295]),
        .I1(out[231]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1311]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1567]_i_16 
       (.I0(\f_permutation_l_/out_reg_n_0_[671] ),
        .I1(\f_permutation_l_/out_reg_n_0_[991] ),
        .I2(\f_permutation_l_/out_reg_n_0_[31] ),
        .I3(\f_permutation_l_/out_reg_n_0_[351] ),
        .O(\out[1567]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1567]_i_17 
       (.I0(\f_permutation_l_/i_reg_n_0_[10] ),
        .I1(\f_permutation_l_/i_reg_n_0_[18] ),
        .I2(\f_permutation_l_/i_reg_n_0_[4] ),
        .I3(\f_permutation_l_/i_reg_n_0_[19] ),
        .I4(\f_permutation_l_/i_reg_n_0_[5] ),
        .I5(\f_permutation_l_/i_reg_n_0_[9] ),
        .O(\out[1567]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1567]_i_2 
       (.I0(\f_permutation_l_/round_in [1203]),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1587]),
        .I4(\out[1567]_i_9_n_0 ),
        .O(\out[1567]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1567]_i_3 
       (.I0(\out[1567]_i_10_n_0 ),
        .I1(padder_out_1[460]),
        .I2(out[396]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1567]_i_11_n_0 ),
        .I5(\f_permutation_l_/round_in [1395]),
        .O(\out[1567]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1567]_i_4 
       (.I0(\f_permutation_l_/round_in [1567]),
        .I1(\f_permutation_l_/round_in [1502]),
        .I2(\out[1545]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[1567]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \out[1567]_i_5 
       (.I0(\out[1567]_i_17_n_0 ),
        .I1(\f_permutation_l_/p_0_in ),
        .I2(\f_permutation_l_/i_reg_n_0_[2] ),
        .I3(\f_permutation_l_/i_reg_n_0_[11] ),
        .I4(\f_permutation_l_/i_reg_n_0_[21] ),
        .O(\f_permutation_l_/rc [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_6 
       (.I0(padder_out_1[394]),
        .I1(out[330]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1458]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1567]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[818] ),
        .I1(padder_out_1[74]),
        .I2(out[10]),
        .I3(\f_permutation_l_/out_reg_n_0_[178] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[498] ),
        .O(\out[1567]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1567]_i_8 
       (.I0(padder_out_1[523]),
        .I1(out[459]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1587]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1567]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[947] ),
        .I1(padder_out_1[203]),
        .I2(out[139]),
        .I3(\f_permutation_l_/out_reg_n_0_[307] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[627] ),
        .O(\out[1567]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1568]_i_1 
       (.I0(\f_permutation_l_/round_in [1204]),
        .I1(\out[1568]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[821] ),
        .I3(\out[1568]_i_4_n_0 ),
        .I4(\out[1568]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1568]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1568]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[756] ),
        .I1(padder_out_1[12]),
        .I2(\f_permutation_l_/out_reg_n_0_[1076] ),
        .I3(\f_permutation_l_/out_reg_n_0_[116] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[436] ),
        .O(\out[1568]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_11 
       (.I0(padder_out_1[332]),
        .I1(out[268]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1396]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_12 
       (.I0(padder_out_1[536]),
        .I1(out[472]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1568]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_13 
       (.I0(padder_out_1[487]),
        .I1(out[423]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1503]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_14 
       (.I0(padder_out_1[280]),
        .I1(out[216]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1312]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1568]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[672] ),
        .I1(\f_permutation_l_/out_reg_n_0_[992] ),
        .I2(\f_permutation_l_/out_reg_n_0_[32] ),
        .I3(\f_permutation_l_/out_reg_n_0_[352] ),
        .O(\out[1568]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_2 
       (.I0(padder_out_1[140]),
        .I1(out[76]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1204]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1568]_i_3 
       (.I0(\out[1568]_i_6_n_0 ),
        .I1(padder_out_1[524]),
        .I2(out[460]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1568]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1459]),
        .O(\out[1568]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1568]_i_4 
       (.I0(\out[1568]_i_9_n_0 ),
        .I1(padder_out_1[461]),
        .I2(out[397]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1568]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1396]),
        .O(\out[1568]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1568]_i_5 
       (.I0(\f_permutation_l_/round_in [1568]),
        .I1(\f_permutation_l_/round_in [1503]),
        .I2(\out[1546]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[1568]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1568]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[948] ),
        .I1(padder_out_1[204]),
        .I2(out[140]),
        .I3(\f_permutation_l_/out_reg_n_0_[308] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[628] ),
        .O(\out[1568]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1568]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[819] ),
        .I1(padder_out_1[75]),
        .I2(out[11]),
        .I3(\f_permutation_l_/out_reg_n_0_[179] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[499] ),
        .O(\out[1568]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1568]_i_8 
       (.I0(padder_out_1[395]),
        .I1(out[331]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1459]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1568]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[885] ),
        .I1(padder_out_1[141]),
        .I2(out[77]),
        .I3(\f_permutation_l_/out_reg_n_0_[245] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[565] ),
        .O(\out[1568]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1569]_i_1 
       (.I0(\f_permutation_l_/round_in [1205]),
        .I1(\out[1569]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[822] ),
        .I3(\out[1569]_i_4_n_0 ),
        .I4(\out[1569]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1569]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1569]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[757] ),
        .I1(padder_out_1[13]),
        .I2(\f_permutation_l_/out_reg_n_0_[1077] ),
        .I3(\f_permutation_l_/out_reg_n_0_[117] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[437] ),
        .O(\out[1569]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_11 
       (.I0(padder_out_1[333]),
        .I1(out[269]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1397]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_12 
       (.I0(padder_out_1[537]),
        .I1(out[473]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1569]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_13 
       (.I0(padder_out_1[472]),
        .I1(out[408]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1504]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_14 
       (.I0(padder_out_1[281]),
        .I1(out[217]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1313]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1569]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[673] ),
        .I1(\f_permutation_l_/out_reg_n_0_[993] ),
        .I2(\f_permutation_l_/out_reg_n_0_[33] ),
        .I3(\f_permutation_l_/out_reg_n_0_[353] ),
        .O(\out[1569]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_2 
       (.I0(padder_out_1[141]),
        .I1(out[77]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1205]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1569]_i_3 
       (.I0(\out[1569]_i_6_n_0 ),
        .I1(padder_out_1[525]),
        .I2(out[461]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1569]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1460]),
        .O(\out[1569]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1569]_i_4 
       (.I0(\out[1569]_i_9_n_0 ),
        .I1(padder_out_1[462]),
        .I2(out[398]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1569]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1397]),
        .O(\out[1569]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1569]_i_5 
       (.I0(\f_permutation_l_/round_in [1569]),
        .I1(\f_permutation_l_/round_in [1504]),
        .I2(\out[1547]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[1569]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1569]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[949] ),
        .I1(padder_out_1[205]),
        .I2(out[141]),
        .I3(\f_permutation_l_/out_reg_n_0_[309] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[629] ),
        .O(\out[1569]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1569]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[820] ),
        .I1(padder_out_1[76]),
        .I2(out[12]),
        .I3(\f_permutation_l_/out_reg_n_0_[180] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[500] ),
        .O(\out[1569]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1569]_i_8 
       (.I0(padder_out_1[396]),
        .I1(out[332]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1460]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1569]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[886] ),
        .I1(padder_out_1[142]),
        .I2(out[78]),
        .I3(\f_permutation_l_/out_reg_n_0_[246] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[566] ),
        .O(\out[1569]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[156]_i_1 
       (.I0(\out[1411]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[693] ),
        .I2(\out[156]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[218] ),
        .I4(\out[1542]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [156]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[156]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[627] ),
        .I1(\f_permutation_l_/round_in [1522]),
        .I2(\out[1565]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[156]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1570]_i_1 
       (.I0(\f_permutation_l_/round_in [1206]),
        .I1(\out[1570]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[823] ),
        .I3(\out[1570]_i_4_n_0 ),
        .I4(\out[1570]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1570]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1570]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[758] ),
        .I1(padder_out_1[14]),
        .I2(\f_permutation_l_/out_reg_n_0_[1078] ),
        .I3(\f_permutation_l_/out_reg_n_0_[118] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[438] ),
        .O(\out[1570]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_11 
       (.I0(padder_out_1[334]),
        .I1(out[270]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1398]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_12 
       (.I0(padder_out_1[538]),
        .I1(out[474]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1570]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_13 
       (.I0(padder_out_1[473]),
        .I1(out[409]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1505]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_14 
       (.I0(padder_out_1[282]),
        .I1(out[218]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1314]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1570]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[674] ),
        .I1(\f_permutation_l_/out_reg_n_0_[994] ),
        .I2(\f_permutation_l_/out_reg_n_0_[34] ),
        .I3(\f_permutation_l_/out_reg_n_0_[354] ),
        .O(\out[1570]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_2 
       (.I0(padder_out_1[142]),
        .I1(out[78]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1206]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1570]_i_3 
       (.I0(\out[1570]_i_6_n_0 ),
        .I1(padder_out_1[526]),
        .I2(out[462]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1570]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1461]),
        .O(\out[1570]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1570]_i_4 
       (.I0(\out[1570]_i_9_n_0 ),
        .I1(padder_out_1[463]),
        .I2(out[399]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1570]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1398]),
        .O(\out[1570]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1570]_i_5 
       (.I0(\f_permutation_l_/round_in [1570]),
        .I1(\f_permutation_l_/round_in [1505]),
        .I2(\out[1548]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[1570]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1570]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[950] ),
        .I1(padder_out_1[206]),
        .I2(out[142]),
        .I3(\f_permutation_l_/out_reg_n_0_[310] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[630] ),
        .O(\out[1570]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1570]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[821] ),
        .I1(padder_out_1[77]),
        .I2(out[13]),
        .I3(\f_permutation_l_/out_reg_n_0_[181] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[501] ),
        .O(\out[1570]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1570]_i_8 
       (.I0(padder_out_1[397]),
        .I1(out[333]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1461]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1570]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[887] ),
        .I1(padder_out_1[143]),
        .I2(out[79]),
        .I3(\f_permutation_l_/out_reg_n_0_[247] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[567] ),
        .O(\out[1570]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1571]_i_1 
       (.I0(\f_permutation_l_/round_in [1207]),
        .I1(\out[1571]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[824] ),
        .I3(\out[1571]_i_4_n_0 ),
        .I4(\out[1571]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1571]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1571]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[759] ),
        .I1(padder_out_1[15]),
        .I2(\f_permutation_l_/out_reg_n_0_[1079] ),
        .I3(\f_permutation_l_/out_reg_n_0_[119] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[439] ),
        .O(\out[1571]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1571]_i_11 
       (.I0(padder_out_1[335]),
        .I1(out[271]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1399]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1571]_i_12 
       (.I0(padder_out_1[474]),
        .I1(out[410]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1506]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1571]_i_13 
       (.I0(padder_out_1[283]),
        .I1(out[219]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1315]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1571]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[675] ),
        .I1(\f_permutation_l_/out_reg_n_0_[995] ),
        .I2(\f_permutation_l_/out_reg_n_0_[35] ),
        .I3(\f_permutation_l_/out_reg_n_0_[355] ),
        .O(\out[1571]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1571]_i_2 
       (.I0(padder_out_1[143]),
        .I1(out[79]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1207]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1571]_i_3 
       (.I0(\out[1571]_i_6_n_0 ),
        .I1(padder_out_1[527]),
        .I2(out[463]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1571]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1462]),
        .O(\out[1571]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1571]_i_4 
       (.I0(\out[1571]_i_9_n_0 ),
        .I1(padder_out_1[448]),
        .I2(out[384]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1571]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1399]),
        .O(\out[1571]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1571]_i_5 
       (.I0(\f_permutation_l_/round_in [1571]),
        .I1(\f_permutation_l_/round_in [1506]),
        .I2(\out[1549]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[1571]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1571]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[951] ),
        .I1(padder_out_1[207]),
        .I2(out[143]),
        .I3(\f_permutation_l_/out_reg_n_0_[311] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[631] ),
        .O(\out[1571]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1571]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[822] ),
        .I1(padder_out_1[78]),
        .I2(out[14]),
        .I3(\f_permutation_l_/out_reg_n_0_[182] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[502] ),
        .O(\out[1571]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1571]_i_8 
       (.I0(padder_out_1[398]),
        .I1(out[334]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1462]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1571]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[888] ),
        .I1(padder_out_1[128]),
        .I2(out[64]),
        .I3(\f_permutation_l_/out_reg_n_0_[248] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[568] ),
        .O(\out[1571]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1572]_i_1 
       (.I0(\f_permutation_l_/round_in [1208]),
        .I1(\out[1572]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[825] ),
        .I3(\out[1572]_i_4_n_0 ),
        .I4(\out[1572]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1572]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1572]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[760] ),
        .I1(padder_out_1[0]),
        .I2(\f_permutation_l_/out_reg_n_0_[1080] ),
        .I3(\f_permutation_l_/out_reg_n_0_[120] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[440] ),
        .O(\out[1572]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_11 
       (.I0(padder_out_1[320]),
        .I1(out[256]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1400]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_12 
       (.I0(padder_out_1[540]),
        .I1(out[476]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1572]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_13 
       (.I0(padder_out_1[475]),
        .I1(out[411]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1507]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_14 
       (.I0(padder_out_1[284]),
        .I1(out[220]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1316]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1572]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[676] ),
        .I1(\f_permutation_l_/out_reg_n_0_[996] ),
        .I2(\f_permutation_l_/out_reg_n_0_[36] ),
        .I3(\f_permutation_l_/out_reg_n_0_[356] ),
        .O(\out[1572]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_2 
       (.I0(padder_out_1[128]),
        .I1(out[64]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1208]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1572]_i_3 
       (.I0(\out[1572]_i_6_n_0 ),
        .I1(padder_out_1[512]),
        .I2(out[448]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1572]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1463]),
        .O(\out[1572]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1572]_i_4 
       (.I0(\out[1572]_i_9_n_0 ),
        .I1(padder_out_1[449]),
        .I2(out[385]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1572]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1400]),
        .O(\out[1572]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1572]_i_5 
       (.I0(\f_permutation_l_/round_in [1572]),
        .I1(\f_permutation_l_/round_in [1507]),
        .I2(\out[1550]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[1572]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1572]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[952] ),
        .I1(padder_out_1[192]),
        .I2(out[128]),
        .I3(\f_permutation_l_/out_reg_n_0_[312] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[632] ),
        .O(\out[1572]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1572]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[823] ),
        .I1(padder_out_1[79]),
        .I2(out[15]),
        .I3(\f_permutation_l_/out_reg_n_0_[183] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[503] ),
        .O(\out[1572]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1572]_i_8 
       (.I0(padder_out_1[399]),
        .I1(out[335]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1463]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1572]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[889] ),
        .I1(padder_out_1[129]),
        .I2(out[65]),
        .I3(\f_permutation_l_/out_reg_n_0_[249] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[569] ),
        .O(\out[1572]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1573]_i_1 
       (.I0(\f_permutation_l_/round_in [1209]),
        .I1(\out[1573]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[826] ),
        .I3(\out[1573]_i_4_n_0 ),
        .I4(\out[1573]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1573]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1573]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[761] ),
        .I1(padder_out_1[1]),
        .I2(\f_permutation_l_/out_reg_n_0_[1081] ),
        .I3(\f_permutation_l_/out_reg_n_0_[121] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[441] ),
        .O(\out[1573]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_11 
       (.I0(padder_out_1[321]),
        .I1(out[257]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1401]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_12 
       (.I0(padder_out_1[541]),
        .I1(out[477]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1573]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_13 
       (.I0(padder_out_1[476]),
        .I1(out[412]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1508]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_14 
       (.I0(padder_out_1[285]),
        .I1(out[221]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1317]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1573]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[677] ),
        .I1(\f_permutation_l_/out_reg_n_0_[997] ),
        .I2(\f_permutation_l_/out_reg_n_0_[37] ),
        .I3(\f_permutation_l_/out_reg_n_0_[357] ),
        .O(\out[1573]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_2 
       (.I0(padder_out_1[129]),
        .I1(out[65]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1209]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1573]_i_3 
       (.I0(\out[1573]_i_6_n_0 ),
        .I1(padder_out_1[513]),
        .I2(out[449]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1573]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1464]),
        .O(\out[1573]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1573]_i_4 
       (.I0(\out[1573]_i_9_n_0 ),
        .I1(padder_out_1[450]),
        .I2(out[386]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1573]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1401]),
        .O(\out[1573]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1573]_i_5 
       (.I0(\f_permutation_l_/round_in [1573]),
        .I1(\f_permutation_l_/round_in [1508]),
        .I2(\out[1551]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[1573]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1573]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[953] ),
        .I1(padder_out_1[193]),
        .I2(out[129]),
        .I3(\f_permutation_l_/out_reg_n_0_[313] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[633] ),
        .O(\out[1573]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1573]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[824] ),
        .I1(padder_out_1[64]),
        .I2(out[0]),
        .I3(\f_permutation_l_/out_reg_n_0_[184] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[504] ),
        .O(\out[1573]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1573]_i_8 
       (.I0(padder_out_1[384]),
        .I1(out[320]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1464]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1573]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[890] ),
        .I1(padder_out_1[130]),
        .I2(out[66]),
        .I3(\f_permutation_l_/out_reg_n_0_[250] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[570] ),
        .O(\out[1573]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1574]_i_1 
       (.I0(\f_permutation_l_/round_in [1210]),
        .I1(\out[1574]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[827] ),
        .I3(\out[1574]_i_4_n_0 ),
        .I4(\out[1574]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1574]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1574]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[762] ),
        .I1(padder_out_1[2]),
        .I2(\f_permutation_l_/out_reg_n_0_[1082] ),
        .I3(\f_permutation_l_/out_reg_n_0_[122] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[442] ),
        .O(\out[1574]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_11 
       (.I0(padder_out_1[322]),
        .I1(out[258]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1402]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_12 
       (.I0(padder_out_1[542]),
        .I1(out[478]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1574]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_13 
       (.I0(padder_out_1[477]),
        .I1(out[413]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1509]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_14 
       (.I0(padder_out_1[286]),
        .I1(out[222]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1318]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1574]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[678] ),
        .I1(\f_permutation_l_/out_reg_n_0_[998] ),
        .I2(\f_permutation_l_/out_reg_n_0_[38] ),
        .I3(\f_permutation_l_/out_reg_n_0_[358] ),
        .O(\out[1574]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_2 
       (.I0(padder_out_1[130]),
        .I1(out[66]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1210]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1574]_i_3 
       (.I0(\out[1574]_i_6_n_0 ),
        .I1(padder_out_1[514]),
        .I2(out[450]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1574]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1465]),
        .O(\out[1574]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1574]_i_4 
       (.I0(\out[1574]_i_9_n_0 ),
        .I1(padder_out_1[451]),
        .I2(out[387]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1574]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1402]),
        .O(\out[1574]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1574]_i_5 
       (.I0(\f_permutation_l_/round_in [1574]),
        .I1(\f_permutation_l_/round_in [1509]),
        .I2(\out[1552]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[1574]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1574]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[954] ),
        .I1(padder_out_1[194]),
        .I2(out[130]),
        .I3(\f_permutation_l_/out_reg_n_0_[314] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[634] ),
        .O(\out[1574]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1574]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[825] ),
        .I1(padder_out_1[65]),
        .I2(out[1]),
        .I3(\f_permutation_l_/out_reg_n_0_[185] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[505] ),
        .O(\out[1574]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1574]_i_8 
       (.I0(padder_out_1[385]),
        .I1(out[321]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1465]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1574]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[891] ),
        .I1(padder_out_1[131]),
        .I2(out[67]),
        .I3(\f_permutation_l_/out_reg_n_0_[251] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[571] ),
        .O(\out[1574]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1575]_i_1 
       (.I0(\f_permutation_l_/round_in [1211]),
        .I1(\out[1575]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[828] ),
        .I3(\out[1575]_i_4_n_0 ),
        .I4(\out[1575]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1575]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1575]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[763] ),
        .I1(padder_out_1[3]),
        .I2(\f_permutation_l_/out_reg_n_0_[1083] ),
        .I3(\f_permutation_l_/out_reg_n_0_[123] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[443] ),
        .O(\out[1575]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_11 
       (.I0(padder_out_1[323]),
        .I1(out[259]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1403]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_12 
       (.I0(padder_out_1[543]),
        .I1(out[479]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1575]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_13 
       (.I0(padder_out_1[478]),
        .I1(out[414]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1510]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_14 
       (.I0(padder_out_1[287]),
        .I1(out[223]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1319]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1575]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[679] ),
        .I1(\f_permutation_l_/out_reg_n_0_[999] ),
        .I2(\f_permutation_l_/out_reg_n_0_[39] ),
        .I3(\f_permutation_l_/out_reg_n_0_[359] ),
        .O(\out[1575]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_2 
       (.I0(padder_out_1[131]),
        .I1(out[67]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1211]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1575]_i_3 
       (.I0(\out[1575]_i_6_n_0 ),
        .I1(padder_out_1[515]),
        .I2(out[451]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1575]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1466]),
        .O(\out[1575]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1575]_i_4 
       (.I0(\out[1575]_i_9_n_0 ),
        .I1(padder_out_1[452]),
        .I2(out[388]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1575]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1403]),
        .O(\out[1575]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1575]_i_5 
       (.I0(\f_permutation_l_/round_in [1575]),
        .I1(\f_permutation_l_/round_in [1510]),
        .I2(\out[1553]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[1575]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1575]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[955] ),
        .I1(padder_out_1[195]),
        .I2(out[131]),
        .I3(\f_permutation_l_/out_reg_n_0_[315] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[635] ),
        .O(\out[1575]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1575]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[826] ),
        .I1(padder_out_1[66]),
        .I2(out[2]),
        .I3(\f_permutation_l_/out_reg_n_0_[186] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[506] ),
        .O(\out[1575]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1575]_i_8 
       (.I0(padder_out_1[386]),
        .I1(out[322]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1466]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1575]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[892] ),
        .I1(padder_out_1[132]),
        .I2(out[68]),
        .I3(\f_permutation_l_/out_reg_n_0_[252] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[572] ),
        .O(\out[1575]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1576]_i_1 
       (.I0(\f_permutation_l_/round_in [1212]),
        .I1(\out[1576]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[829] ),
        .I3(\out[1576]_i_4_n_0 ),
        .I4(\out[1576]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1576]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1576]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[764] ),
        .I1(padder_out_1[4]),
        .I2(\f_permutation_l_/out_reg_n_0_[1084] ),
        .I3(\f_permutation_l_/out_reg_n_0_[124] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[444] ),
        .O(\out[1576]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_11 
       (.I0(padder_out_1[324]),
        .I1(out[260]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1404]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_12 
       (.I0(padder_out_1[528]),
        .I1(out[464]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1576]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_13 
       (.I0(padder_out_1[479]),
        .I1(out[415]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1511]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_14 
       (.I0(padder_out_1[272]),
        .I1(out[208]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1320]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1576]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[680] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1000] ),
        .I2(\f_permutation_l_/out_reg_n_0_[40] ),
        .I3(\f_permutation_l_/out_reg_n_0_[360] ),
        .O(\out[1576]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_2 
       (.I0(padder_out_1[132]),
        .I1(out[68]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1212]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1576]_i_3 
       (.I0(\out[1576]_i_6_n_0 ),
        .I1(padder_out_1[516]),
        .I2(out[452]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1576]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1467]),
        .O(\out[1576]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1576]_i_4 
       (.I0(\out[1576]_i_9_n_0 ),
        .I1(padder_out_1[453]),
        .I2(out[389]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1576]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1404]),
        .O(\out[1576]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1576]_i_5 
       (.I0(\f_permutation_l_/round_in [1576]),
        .I1(\f_permutation_l_/round_in [1511]),
        .I2(\out[1554]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[1576]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1576]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[956] ),
        .I1(padder_out_1[196]),
        .I2(out[132]),
        .I3(\f_permutation_l_/out_reg_n_0_[316] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[636] ),
        .O(\out[1576]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1576]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[827] ),
        .I1(padder_out_1[67]),
        .I2(out[3]),
        .I3(\f_permutation_l_/out_reg_n_0_[187] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[507] ),
        .O(\out[1576]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1576]_i_8 
       (.I0(padder_out_1[387]),
        .I1(out[323]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1467]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1576]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[893] ),
        .I1(padder_out_1[133]),
        .I2(out[69]),
        .I3(\f_permutation_l_/out_reg_n_0_[253] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[573] ),
        .O(\out[1576]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[1577]_i_1 
       (.I0(\f_permutation_l_/round_in [1213]),
        .I1(\out[1577]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[830] ),
        .I3(\out[1577]_i_4_n_0 ),
        .I4(\out[1577]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1577]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1577]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[765] ),
        .I1(padder_out_1[5]),
        .I2(\f_permutation_l_/out_reg_n_0_[1085] ),
        .I3(\f_permutation_l_/out_reg_n_0_[125] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[445] ),
        .O(\out[1577]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_11 
       (.I0(padder_out_1[325]),
        .I1(out[261]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1405]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_12 
       (.I0(padder_out_1[529]),
        .I1(out[465]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1577]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_13 
       (.I0(padder_out_1[464]),
        .I1(out[400]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1512]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_14 
       (.I0(padder_out_1[273]),
        .I1(out[209]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1321]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1577]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[681] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1001] ),
        .I2(\f_permutation_l_/out_reg_n_0_[41] ),
        .I3(\f_permutation_l_/out_reg_n_0_[361] ),
        .O(\out[1577]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_2 
       (.I0(padder_out_1[133]),
        .I1(out[69]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1213]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1577]_i_3 
       (.I0(\out[1577]_i_6_n_0 ),
        .I1(padder_out_1[517]),
        .I2(out[453]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1577]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1468]),
        .O(\out[1577]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1577]_i_4 
       (.I0(\out[1577]_i_9_n_0 ),
        .I1(padder_out_1[454]),
        .I2(out[390]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1577]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1405]),
        .O(\out[1577]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1577]_i_5 
       (.I0(\f_permutation_l_/round_in [1577]),
        .I1(\f_permutation_l_/round_in [1512]),
        .I2(\out[1555]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[1577]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1577]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[957] ),
        .I1(padder_out_1[197]),
        .I2(out[133]),
        .I3(\f_permutation_l_/out_reg_n_0_[317] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[637] ),
        .O(\out[1577]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1577]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[828] ),
        .I1(padder_out_1[68]),
        .I2(out[4]),
        .I3(\f_permutation_l_/out_reg_n_0_[188] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[508] ),
        .O(\out[1577]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1577]_i_8 
       (.I0(padder_out_1[388]),
        .I1(out[324]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1468]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1577]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[894] ),
        .I1(padder_out_1[134]),
        .I2(out[70]),
        .I3(\f_permutation_l_/out_reg_n_0_[254] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[574] ),
        .O(\out[1577]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1578]_i_1 
       (.I0(\f_permutation_l_/round_in [1214]),
        .I1(\out[1578]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[831] ),
        .I3(\out[1578]_i_4_n_0 ),
        .I4(\out[1578]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1578]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_10 
       (.I0(padder_out_1[326]),
        .I1(out[262]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1406]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_11 
       (.I0(padder_out_1[530]),
        .I1(out[466]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1578]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_12 
       (.I0(padder_out_1[465]),
        .I1(out[401]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1513]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_13 
       (.I0(padder_out_1[274]),
        .I1(out[210]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1322]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1578]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[682] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1002] ),
        .I2(\f_permutation_l_/out_reg_n_0_[42] ),
        .I3(\f_permutation_l_/out_reg_n_0_[362] ),
        .O(\out[1578]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_2 
       (.I0(padder_out_1[134]),
        .I1(out[70]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1214]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1578]_i_3 
       (.I0(\out[1578]_i_6_n_0 ),
        .I1(padder_out_1[518]),
        .I2(out[454]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1578]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1469]),
        .O(\out[1578]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1578]_i_4 
       (.I0(\out[1536]_i_19_n_0 ),
        .I1(padder_out_1[455]),
        .I2(out[391]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1578]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1406]),
        .O(\out[1578]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1578]_i_5 
       (.I0(\f_permutation_l_/round_in [1578]),
        .I1(\f_permutation_l_/round_in [1513]),
        .I2(\out[1556]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[1578]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1578]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[958] ),
        .I1(padder_out_1[198]),
        .I2(out[134]),
        .I3(\f_permutation_l_/out_reg_n_0_[318] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[638] ),
        .O(\out[1578]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1578]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[829] ),
        .I1(padder_out_1[69]),
        .I2(out[5]),
        .I3(\f_permutation_l_/out_reg_n_0_[189] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[509] ),
        .O(\out[1578]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1578]_i_8 
       (.I0(padder_out_1[389]),
        .I1(out[325]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1469]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1578]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[766] ),
        .I1(padder_out_1[6]),
        .I2(\f_permutation_l_/out_reg_n_0_[1086] ),
        .I3(\f_permutation_l_/out_reg_n_0_[126] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[446] ),
        .O(\out[1578]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1579]_i_1 
       (.I0(\f_permutation_l_/round_in [1215]),
        .I1(\out[1579]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[768] ),
        .I3(\out[1579]_i_4_n_0 ),
        .I4(\out[1579]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1579]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1579]_i_10 
       (.I0(\f_permutation_l_/out_reg_n_0_[767] ),
        .I1(padder_out_1[7]),
        .I2(\f_permutation_l_/out_reg_n_0_[1087] ),
        .I3(\f_permutation_l_/out_reg_n_0_[127] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[447] ),
        .O(\out[1579]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_11 
       (.I0(padder_out_1[327]),
        .I1(out[263]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1407]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_12 
       (.I0(padder_out_1[531]),
        .I1(out[467]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1579]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_13 
       (.I0(padder_out_1[466]),
        .I1(out[402]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1514]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_14 
       (.I0(padder_out_1[275]),
        .I1(out[211]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1323]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1579]_i_15 
       (.I0(\f_permutation_l_/out_reg_n_0_[683] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1003] ),
        .I2(\f_permutation_l_/out_reg_n_0_[43] ),
        .I3(\f_permutation_l_/out_reg_n_0_[363] ),
        .O(\out[1579]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_2 
       (.I0(padder_out_1[135]),
        .I1(out[71]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1215]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1579]_i_3 
       (.I0(\out[1579]_i_7_n_0 ),
        .I1(padder_out_1[519]),
        .I2(out[455]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1579]_i_8_n_0 ),
        .I5(\f_permutation_l_/round_in [1470]),
        .O(\out[1579]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1579]_i_4 
       (.I0(\out[1537]_i_17_n_0 ),
        .I1(padder_out_1[504]),
        .I2(out[440]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1579]_i_10_n_0 ),
        .I5(\f_permutation_l_/round_in [1407]),
        .O(\out[1579]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1579]_i_5 
       (.I0(\f_permutation_l_/round_in [1579]),
        .I1(\f_permutation_l_/round_in [1514]),
        .I2(\out[1557]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[1579]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[1579]_i_6 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[1579]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1579]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[959] ),
        .I1(padder_out_1[199]),
        .I2(out[135]),
        .I3(\f_permutation_l_/out_reg_n_0_[319] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[639] ),
        .O(\out[1579]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1579]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[830] ),
        .I1(padder_out_1[70]),
        .I2(out[6]),
        .I3(\f_permutation_l_/out_reg_n_0_[190] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[510] ),
        .O(\out[1579]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1579]_i_9 
       (.I0(padder_out_1[390]),
        .I1(out[326]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1470]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[157]_i_1 
       (.I0(\out[1412]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[694] ),
        .I2(\out[157]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[219] ),
        .I4(\out[1287]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [157]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[157]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[628] ),
        .I1(\f_permutation_l_/round_in [1523]),
        .I2(\out[1566]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[157]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1580]_i_1 
       (.I0(\f_permutation_l_/round_in [1152]),
        .I1(\out[1580]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[769] ),
        .I3(\out[1580]_i_4_n_0 ),
        .I4(\out[1580]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1580]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_10 
       (.I0(padder_out_1[376]),
        .I1(out[312]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1344]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_11 
       (.I0(padder_out_1[532]),
        .I1(out[468]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1580]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_12 
       (.I0(padder_out_1[467]),
        .I1(out[403]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1515]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_13 
       (.I0(padder_out_1[276]),
        .I1(out[212]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1324]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1580]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[684] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1004] ),
        .I2(\f_permutation_l_/out_reg_n_0_[44] ),
        .I3(\f_permutation_l_/out_reg_n_0_[364] ),
        .O(\out[1580]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_2 
       (.I0(padder_out_1[184]),
        .I1(out[120]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1152]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1580]_i_3 
       (.I0(\out[1580]_i_6_n_0 ),
        .I1(padder_out_1[568]),
        .I2(out[504]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1580]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1471]),
        .O(\out[1580]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1580]_i_4 
       (.I0(\out[1538]_i_16_n_0 ),
        .I1(padder_out_1[505]),
        .I2(out[441]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1580]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1344]),
        .O(\out[1580]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1580]_i_5 
       (.I0(\f_permutation_l_/round_in [1580]),
        .I1(\f_permutation_l_/round_in [1515]),
        .I2(\out[1558]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[1580]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1580]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[896] ),
        .I1(padder_out_1[248]),
        .I2(out[184]),
        .I3(\f_permutation_l_/out_reg_n_0_[256] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[576] ),
        .O(\out[1580]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1580]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[831] ),
        .I1(padder_out_1[71]),
        .I2(out[7]),
        .I3(\f_permutation_l_/out_reg_n_0_[191] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[511] ),
        .O(\out[1580]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1580]_i_8 
       (.I0(padder_out_1[391]),
        .I1(out[327]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1471]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1580]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[704] ),
        .I1(padder_out_1[56]),
        .I2(\f_permutation_l_/out_reg_n_0_[1024] ),
        .I3(\f_permutation_l_/out_reg_n_0_[64] ),
        .I4(\out[1543]_i_23_n_0 ),
        .I5(\f_permutation_l_/out_reg_n_0_[384] ),
        .O(\out[1580]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[1581]_i_1 
       (.I0(\f_permutation_l_/round_in [1153]),
        .I1(\out[1581]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[770] ),
        .I3(\out[1581]_i_4_n_0 ),
        .I4(\out[1581]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1581]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_10 
       (.I0(padder_out_1[377]),
        .I1(out[313]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1345]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_11 
       (.I0(padder_out_1[533]),
        .I1(out[469]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1581]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_12 
       (.I0(padder_out_1[468]),
        .I1(out[404]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1516]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_13 
       (.I0(padder_out_1[277]),
        .I1(out[213]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1325]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1581]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[685] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1005] ),
        .I2(\f_permutation_l_/out_reg_n_0_[45] ),
        .I3(\f_permutation_l_/out_reg_n_0_[365] ),
        .O(\out[1581]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_2 
       (.I0(padder_out_1[185]),
        .I1(out[121]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1153]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1581]_i_3 
       (.I0(\out[1581]_i_6_n_0 ),
        .I1(padder_out_1[569]),
        .I2(out[505]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1581]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1408]),
        .O(\out[1581]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1581]_i_4 
       (.I0(\out[1539]_i_15_n_0 ),
        .I1(padder_out_1[506]),
        .I2(out[442]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1581]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1345]),
        .O(\out[1581]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1581]_i_5 
       (.I0(\f_permutation_l_/round_in [1581]),
        .I1(\f_permutation_l_/round_in [1516]),
        .I2(\out[1559]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[1581]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1581]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[897] ),
        .I1(padder_out_1[249]),
        .I2(out[185]),
        .I3(\f_permutation_l_/out_reg_n_0_[257] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[577] ),
        .O(\out[1581]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1581]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[768] ),
        .I1(padder_out_1[120]),
        .I2(out[56]),
        .I3(\f_permutation_l_/out_reg_n_0_[128] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[448] ),
        .O(\out[1581]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1581]_i_8 
       (.I0(padder_out_1[440]),
        .I1(out[376]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1408]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1581]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[705] ),
        .I1(padder_out_1[57]),
        .I2(\f_permutation_l_/out_reg_n_0_[1025] ),
        .I3(\f_permutation_l_/out_reg_n_0_[65] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[385] ),
        .O(\out[1581]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1582]_i_1 
       (.I0(\f_permutation_l_/round_in [1154]),
        .I1(\out[1582]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[771] ),
        .I3(\out[1582]_i_4_n_0 ),
        .I4(\out[1582]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1582]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_10 
       (.I0(padder_out_1[378]),
        .I1(out[314]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1346]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_11 
       (.I0(padder_out_1[534]),
        .I1(out[470]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1582]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_12 
       (.I0(padder_out_1[469]),
        .I1(out[405]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1517]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_13 
       (.I0(padder_out_1[278]),
        .I1(out[214]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1326]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1582]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[686] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1006] ),
        .I2(\f_permutation_l_/out_reg_n_0_[46] ),
        .I3(\f_permutation_l_/out_reg_n_0_[366] ),
        .O(\out[1582]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_2 
       (.I0(padder_out_1[186]),
        .I1(out[122]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1154]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1582]_i_3 
       (.I0(\out[1582]_i_6_n_0 ),
        .I1(padder_out_1[570]),
        .I2(out[506]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1582]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1409]),
        .O(\out[1582]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1582]_i_4 
       (.I0(\out[1540]_i_16_n_0 ),
        .I1(padder_out_1[507]),
        .I2(out[443]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1582]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1346]),
        .O(\out[1582]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1582]_i_5 
       (.I0(\f_permutation_l_/round_in [1582]),
        .I1(\f_permutation_l_/round_in [1517]),
        .I2(\out[1560]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[1582]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1582]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[898] ),
        .I1(padder_out_1[250]),
        .I2(out[186]),
        .I3(\f_permutation_l_/out_reg_n_0_[258] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[578] ),
        .O(\out[1582]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1582]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[769] ),
        .I1(padder_out_1[121]),
        .I2(out[57]),
        .I3(\f_permutation_l_/out_reg_n_0_[129] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[449] ),
        .O(\out[1582]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1582]_i_8 
       (.I0(padder_out_1[441]),
        .I1(out[377]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1409]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1582]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[706] ),
        .I1(padder_out_1[58]),
        .I2(\f_permutation_l_/out_reg_n_0_[1026] ),
        .I3(\f_permutation_l_/out_reg_n_0_[66] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[386] ),
        .O(\out[1582]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1583]_i_1 
       (.I0(\f_permutation_l_/round_in [1155]),
        .I1(\out[1583]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[772] ),
        .I3(\out[1583]_i_4_n_0 ),
        .I4(\out[1583]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1583]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_10 
       (.I0(padder_out_1[379]),
        .I1(out[315]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1347]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_11 
       (.I0(padder_out_1[535]),
        .I1(out[471]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1583]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_12 
       (.I0(padder_out_1[470]),
        .I1(out[406]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1518]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_13 
       (.I0(padder_out_1[279]),
        .I1(out[215]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1327]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1583]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[687] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1007] ),
        .I2(\f_permutation_l_/out_reg_n_0_[47] ),
        .I3(\f_permutation_l_/out_reg_n_0_[367] ),
        .O(\out[1583]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_2 
       (.I0(padder_out_1[187]),
        .I1(out[123]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1155]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1583]_i_3 
       (.I0(\out[1583]_i_6_n_0 ),
        .I1(padder_out_1[571]),
        .I2(out[507]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1583]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1410]),
        .O(\out[1583]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1583]_i_4 
       (.I0(\out[1541]_i_16_n_0 ),
        .I1(padder_out_1[508]),
        .I2(out[444]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1583]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1347]),
        .O(\out[1583]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1583]_i_5 
       (.I0(\f_permutation_l_/round_in [1583]),
        .I1(\f_permutation_l_/round_in [1518]),
        .I2(\out[1561]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[1583]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1583]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[899] ),
        .I1(padder_out_1[251]),
        .I2(out[187]),
        .I3(\f_permutation_l_/out_reg_n_0_[259] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[579] ),
        .O(\out[1583]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1583]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[770] ),
        .I1(padder_out_1[122]),
        .I2(out[58]),
        .I3(\f_permutation_l_/out_reg_n_0_[130] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[450] ),
        .O(\out[1583]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1583]_i_8 
       (.I0(padder_out_1[442]),
        .I1(out[378]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1410]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1583]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[707] ),
        .I1(padder_out_1[59]),
        .I2(\f_permutation_l_/out_reg_n_0_[1027] ),
        .I3(\f_permutation_l_/out_reg_n_0_[67] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[387] ),
        .O(\out[1583]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1584]_i_1 
       (.I0(\f_permutation_l_/round_in [1156]),
        .I1(\out[1584]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[773] ),
        .I3(\out[1584]_i_4_n_0 ),
        .I4(\out[1584]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1584]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_10 
       (.I0(padder_out_1[380]),
        .I1(out[316]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1348]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_11 
       (.I0(padder_out_1[520]),
        .I1(out[456]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1584]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_12 
       (.I0(padder_out_1[471]),
        .I1(out[407]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1519]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_13 
       (.I0(padder_out_1[264]),
        .I1(out[200]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1328]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1584]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[688] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1008] ),
        .I2(\f_permutation_l_/out_reg_n_0_[48] ),
        .I3(\f_permutation_l_/out_reg_n_0_[368] ),
        .O(\out[1584]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_2 
       (.I0(padder_out_1[188]),
        .I1(out[124]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1156]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1584]_i_3 
       (.I0(\out[1584]_i_6_n_0 ),
        .I1(padder_out_1[572]),
        .I2(out[508]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1584]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1411]),
        .O(\out[1584]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1584]_i_4 
       (.I0(\out[1542]_i_18_n_0 ),
        .I1(padder_out_1[509]),
        .I2(out[445]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1584]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1348]),
        .O(\out[1584]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1584]_i_5 
       (.I0(\f_permutation_l_/round_in [1584]),
        .I1(\f_permutation_l_/round_in [1519]),
        .I2(\out[1562]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[1584]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1584]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[900] ),
        .I1(padder_out_1[252]),
        .I2(out[188]),
        .I3(\f_permutation_l_/out_reg_n_0_[260] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[580] ),
        .O(\out[1584]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1584]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[771] ),
        .I1(padder_out_1[123]),
        .I2(out[59]),
        .I3(\f_permutation_l_/out_reg_n_0_[131] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[451] ),
        .O(\out[1584]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1584]_i_8 
       (.I0(padder_out_1[443]),
        .I1(out[379]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1411]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1584]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[708] ),
        .I1(padder_out_1[60]),
        .I2(\f_permutation_l_/out_reg_n_0_[1028] ),
        .I3(\f_permutation_l_/out_reg_n_0_[68] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[388] ),
        .O(\out[1584]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1585]_i_1 
       (.I0(\f_permutation_l_/round_in [1157]),
        .I1(\out[1585]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[774] ),
        .I3(\out[1585]_i_4_n_0 ),
        .I4(\out[1585]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1585]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_10 
       (.I0(padder_out_1[381]),
        .I1(out[317]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1349]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_11 
       (.I0(padder_out_1[521]),
        .I1(out[457]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1585]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_12 
       (.I0(padder_out_1[456]),
        .I1(out[392]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1520]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_13 
       (.I0(padder_out_1[265]),
        .I1(out[201]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1329]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1585]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[689] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1009] ),
        .I2(\f_permutation_l_/out_reg_n_0_[49] ),
        .I3(\f_permutation_l_/out_reg_n_0_[369] ),
        .O(\out[1585]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_2 
       (.I0(padder_out_1[189]),
        .I1(out[125]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1157]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1585]_i_3 
       (.I0(\out[1585]_i_6_n_0 ),
        .I1(padder_out_1[573]),
        .I2(out[509]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1585]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1412]),
        .O(\out[1585]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1585]_i_4 
       (.I0(\out[1543]_i_19_n_0 ),
        .I1(padder_out_1[510]),
        .I2(out[446]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1585]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1349]),
        .O(\out[1585]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1585]_i_5 
       (.I0(\f_permutation_l_/round_in [1585]),
        .I1(\f_permutation_l_/round_in [1520]),
        .I2(\out[1563]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[1585]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1585]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[901] ),
        .I1(padder_out_1[253]),
        .I2(out[189]),
        .I3(\f_permutation_l_/out_reg_n_0_[261] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[581] ),
        .O(\out[1585]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1585]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[772] ),
        .I1(padder_out_1[124]),
        .I2(out[60]),
        .I3(\f_permutation_l_/out_reg_n_0_[132] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[452] ),
        .O(\out[1585]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1585]_i_8 
       (.I0(padder_out_1[444]),
        .I1(out[380]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1412]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1585]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[709] ),
        .I1(padder_out_1[61]),
        .I2(\f_permutation_l_/out_reg_n_0_[1029] ),
        .I3(\f_permutation_l_/out_reg_n_0_[69] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[389] ),
        .O(\out[1585]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1586]_i_1 
       (.I0(\f_permutation_l_/round_in [1158]),
        .I1(\out[1586]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[775] ),
        .I3(\out[1586]_i_4_n_0 ),
        .I4(\out[1586]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1586]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_10 
       (.I0(padder_out_1[382]),
        .I1(out[318]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1350]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_11 
       (.I0(padder_out_1[522]),
        .I1(out[458]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1586]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_12 
       (.I0(padder_out_1[457]),
        .I1(out[393]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1521]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_13 
       (.I0(padder_out_1[266]),
        .I1(out[202]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1330]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1586]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[690] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1010] ),
        .I2(\f_permutation_l_/out_reg_n_0_[50] ),
        .I3(\f_permutation_l_/out_reg_n_0_[370] ),
        .O(\out[1586]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_2 
       (.I0(padder_out_1[190]),
        .I1(out[126]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1158]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1586]_i_3 
       (.I0(\out[1586]_i_6_n_0 ),
        .I1(padder_out_1[574]),
        .I2(out[510]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1586]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1413]),
        .O(\out[1586]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1586]_i_4 
       (.I0(\out[1544]_i_16_n_0 ),
        .I1(padder_out_1[511]),
        .I2(out[447]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1586]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1350]),
        .O(\out[1586]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1586]_i_5 
       (.I0(\f_permutation_l_/round_in [1586]),
        .I1(\f_permutation_l_/round_in [1521]),
        .I2(\out[1564]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[1586]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1586]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[902] ),
        .I1(padder_out_1[254]),
        .I2(out[190]),
        .I3(\f_permutation_l_/out_reg_n_0_[262] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[582] ),
        .O(\out[1586]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1586]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[773] ),
        .I1(padder_out_1[125]),
        .I2(out[61]),
        .I3(\f_permutation_l_/out_reg_n_0_[133] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[453] ),
        .O(\out[1586]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1586]_i_8 
       (.I0(padder_out_1[445]),
        .I1(out[381]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1413]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1586]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[710] ),
        .I1(padder_out_1[62]),
        .I2(\f_permutation_l_/out_reg_n_0_[1030] ),
        .I3(\f_permutation_l_/out_reg_n_0_[70] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[390] ),
        .O(\out[1586]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1587]_i_1 
       (.I0(\f_permutation_l_/round_in [1159]),
        .I1(\out[1587]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[776] ),
        .I3(\out[1587]_i_4_n_0 ),
        .I4(\out[1587]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1587]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1587]_i_10 
       (.I0(padder_out_1[383]),
        .I1(out[319]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1351]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1587]_i_11 
       (.I0(padder_out_1[458]),
        .I1(out[394]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1522]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1587]_i_12 
       (.I0(padder_out_1[267]),
        .I1(out[203]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1331]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1587]_i_13 
       (.I0(\f_permutation_l_/out_reg_n_0_[691] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1011] ),
        .I2(\f_permutation_l_/out_reg_n_0_[51] ),
        .I3(\f_permutation_l_/out_reg_n_0_[371] ),
        .O(\out[1587]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1587]_i_2 
       (.I0(padder_out_1[191]),
        .I1(out[127]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1159]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1587]_i_3 
       (.I0(\out[1587]_i_6_n_0 ),
        .I1(padder_out_1[575]),
        .I2(out[511]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1587]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1414]),
        .O(\out[1587]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1587]_i_4 
       (.I0(\out[1545]_i_16_n_0 ),
        .I1(padder_out_1[496]),
        .I2(out[432]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1587]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1351]),
        .O(\out[1587]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1587]_i_5 
       (.I0(\f_permutation_l_/round_in [1587]),
        .I1(\f_permutation_l_/round_in [1522]),
        .I2(\out[1565]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[1587]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1587]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[903] ),
        .I1(padder_out_1[255]),
        .I2(out[191]),
        .I3(\f_permutation_l_/out_reg_n_0_[263] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[583] ),
        .O(\out[1587]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1587]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[774] ),
        .I1(padder_out_1[126]),
        .I2(out[62]),
        .I3(\f_permutation_l_/out_reg_n_0_[134] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[454] ),
        .O(\out[1587]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1587]_i_8 
       (.I0(padder_out_1[446]),
        .I1(out[382]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1414]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1587]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[711] ),
        .I1(padder_out_1[63]),
        .I2(\f_permutation_l_/out_reg_n_0_[1031] ),
        .I3(\f_permutation_l_/out_reg_n_0_[71] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[391] ),
        .O(\out[1587]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1588]_i_1 
       (.I0(\f_permutation_l_/round_in [1160]),
        .I1(\out[1588]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[777] ),
        .I3(\out[1588]_i_4_n_0 ),
        .I4(\out[1588]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1588]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_10 
       (.I0(padder_out_1[368]),
        .I1(out[304]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1352]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_11 
       (.I0(padder_out_1[524]),
        .I1(out[460]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1588]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_12 
       (.I0(padder_out_1[459]),
        .I1(out[395]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1523]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_13 
       (.I0(padder_out_1[268]),
        .I1(out[204]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1332]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1588]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[692] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1012] ),
        .I2(\f_permutation_l_/out_reg_n_0_[52] ),
        .I3(\f_permutation_l_/out_reg_n_0_[372] ),
        .O(\out[1588]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_2 
       (.I0(padder_out_1[176]),
        .I1(out[112]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1160]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1588]_i_3 
       (.I0(\out[1588]_i_6_n_0 ),
        .I1(padder_out_1[560]),
        .I2(out[496]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1588]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1415]),
        .O(\out[1588]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1588]_i_4 
       (.I0(\out[1546]_i_16_n_0 ),
        .I1(padder_out_1[497]),
        .I2(out[433]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1588]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1352]),
        .O(\out[1588]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1588]_i_5 
       (.I0(\f_permutation_l_/round_in [1588]),
        .I1(\f_permutation_l_/round_in [1523]),
        .I2(\out[1566]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[1588]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1588]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[904] ),
        .I1(padder_out_1[240]),
        .I2(out[176]),
        .I3(\f_permutation_l_/out_reg_n_0_[264] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[584] ),
        .O(\out[1588]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1588]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[775] ),
        .I1(padder_out_1[127]),
        .I2(out[63]),
        .I3(\f_permutation_l_/out_reg_n_0_[135] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[455] ),
        .O(\out[1588]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1588]_i_8 
       (.I0(padder_out_1[447]),
        .I1(out[383]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1415]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1588]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[712] ),
        .I1(padder_out_1[48]),
        .I2(\f_permutation_l_/out_reg_n_0_[1032] ),
        .I3(\f_permutation_l_/out_reg_n_0_[72] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[392] ),
        .O(\out[1588]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1589]_i_1 
       (.I0(\f_permutation_l_/round_in [1161]),
        .I1(\out[1589]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[778] ),
        .I3(\out[1589]_i_4_n_0 ),
        .I4(\out[1589]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1589]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_10 
       (.I0(padder_out_1[369]),
        .I1(out[305]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1353]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_11 
       (.I0(padder_out_1[525]),
        .I1(out[461]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1589]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_12 
       (.I0(padder_out_1[460]),
        .I1(out[396]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1524]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_13 
       (.I0(padder_out_1[269]),
        .I1(out[205]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1333]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1589]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[693] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1013] ),
        .I2(\f_permutation_l_/out_reg_n_0_[53] ),
        .I3(\f_permutation_l_/out_reg_n_0_[373] ),
        .O(\out[1589]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_2 
       (.I0(padder_out_1[177]),
        .I1(out[113]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1161]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1589]_i_3 
       (.I0(\out[1589]_i_6_n_0 ),
        .I1(padder_out_1[561]),
        .I2(out[497]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1589]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1416]),
        .O(\out[1589]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1589]_i_4 
       (.I0(\out[1547]_i_16_n_0 ),
        .I1(padder_out_1[498]),
        .I2(out[434]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1589]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1353]),
        .O(\out[1589]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1589]_i_5 
       (.I0(\f_permutation_l_/round_in [1589]),
        .I1(\f_permutation_l_/round_in [1524]),
        .I2(\out[1567]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[1589]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1589]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[905] ),
        .I1(padder_out_1[241]),
        .I2(out[177]),
        .I3(\f_permutation_l_/out_reg_n_0_[265] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[585] ),
        .O(\out[1589]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1589]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[776] ),
        .I1(padder_out_1[112]),
        .I2(out[48]),
        .I3(\f_permutation_l_/out_reg_n_0_[136] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[456] ),
        .O(\out[1589]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1589]_i_8 
       (.I0(padder_out_1[432]),
        .I1(out[368]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1416]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1589]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[713] ),
        .I1(padder_out_1[49]),
        .I2(\f_permutation_l_/out_reg_n_0_[1033] ),
        .I3(\f_permutation_l_/out_reg_n_0_[73] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[393] ),
        .O(\out[1589]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[158]_i_1 
       (.I0(\out[1413]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[695] ),
        .I2(\out[158]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[220] ),
        .I4(\out[1544]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [158]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[158]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[629] ),
        .I1(\f_permutation_l_/round_in [1524]),
        .I2(\out[1567]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[158]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1590]_i_1 
       (.I0(\f_permutation_l_/round_in [1162]),
        .I1(\out[1590]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[779] ),
        .I3(\out[1590]_i_4_n_0 ),
        .I4(\out[1590]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1590]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_10 
       (.I0(padder_out_1[370]),
        .I1(out[306]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1354]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_11 
       (.I0(padder_out_1[526]),
        .I1(out[462]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1590]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_12 
       (.I0(padder_out_1[461]),
        .I1(out[397]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1525]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_13 
       (.I0(padder_out_1[270]),
        .I1(out[206]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1334]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1590]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[694] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1014] ),
        .I2(\f_permutation_l_/out_reg_n_0_[54] ),
        .I3(\f_permutation_l_/out_reg_n_0_[374] ),
        .O(\out[1590]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_2 
       (.I0(padder_out_1[178]),
        .I1(out[114]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1162]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1590]_i_3 
       (.I0(\out[1590]_i_6_n_0 ),
        .I1(padder_out_1[562]),
        .I2(out[498]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1590]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1417]),
        .O(\out[1590]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1590]_i_4 
       (.I0(\out[1548]_i_16_n_0 ),
        .I1(padder_out_1[499]),
        .I2(out[435]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1590]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1354]),
        .O(\out[1590]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1590]_i_5 
       (.I0(\f_permutation_l_/round_in [1590]),
        .I1(\f_permutation_l_/round_in [1525]),
        .I2(\out[1568]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[1590]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1590]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[906] ),
        .I1(padder_out_1[242]),
        .I2(out[178]),
        .I3(\f_permutation_l_/out_reg_n_0_[266] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[586] ),
        .O(\out[1590]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1590]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[777] ),
        .I1(padder_out_1[113]),
        .I2(out[49]),
        .I3(\f_permutation_l_/out_reg_n_0_[137] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[457] ),
        .O(\out[1590]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1590]_i_8 
       (.I0(padder_out_1[433]),
        .I1(out[369]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1417]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1590]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[714] ),
        .I1(padder_out_1[50]),
        .I2(\f_permutation_l_/out_reg_n_0_[1034] ),
        .I3(\f_permutation_l_/out_reg_n_0_[74] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[394] ),
        .O(\out[1590]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1591]_i_1 
       (.I0(\f_permutation_l_/round_in [1163]),
        .I1(\out[1591]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[780] ),
        .I3(\out[1591]_i_4_n_0 ),
        .I4(\out[1591]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1591]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_10 
       (.I0(padder_out_1[371]),
        .I1(out[307]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1355]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_11 
       (.I0(padder_out_1[527]),
        .I1(out[463]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1591]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_12 
       (.I0(padder_out_1[462]),
        .I1(out[398]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1526]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_13 
       (.I0(padder_out_1[271]),
        .I1(out[207]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1335]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1591]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[695] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1015] ),
        .I2(\f_permutation_l_/out_reg_n_0_[55] ),
        .I3(\f_permutation_l_/out_reg_n_0_[375] ),
        .O(\out[1591]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_2 
       (.I0(padder_out_1[179]),
        .I1(out[115]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1163]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1591]_i_3 
       (.I0(\out[1591]_i_6_n_0 ),
        .I1(padder_out_1[563]),
        .I2(out[499]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1591]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1418]),
        .O(\out[1591]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1591]_i_4 
       (.I0(\out[1549]_i_16_n_0 ),
        .I1(padder_out_1[500]),
        .I2(out[436]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1591]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1355]),
        .O(\out[1591]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1591]_i_5 
       (.I0(\f_permutation_l_/round_in [1591]),
        .I1(\f_permutation_l_/round_in [1526]),
        .I2(\out[1569]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[1591]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1591]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[907] ),
        .I1(padder_out_1[243]),
        .I2(out[179]),
        .I3(\f_permutation_l_/out_reg_n_0_[267] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[587] ),
        .O(\out[1591]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1591]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[778] ),
        .I1(padder_out_1[114]),
        .I2(out[50]),
        .I3(\f_permutation_l_/out_reg_n_0_[138] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[458] ),
        .O(\out[1591]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1591]_i_8 
       (.I0(padder_out_1[434]),
        .I1(out[370]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1418]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1591]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[715] ),
        .I1(padder_out_1[51]),
        .I2(\f_permutation_l_/out_reg_n_0_[1035] ),
        .I3(\f_permutation_l_/out_reg_n_0_[75] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[395] ),
        .O(\out[1591]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1592]_i_1 
       (.I0(\f_permutation_l_/round_in [1164]),
        .I1(\out[1592]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[781] ),
        .I3(\out[1592]_i_4_n_0 ),
        .I4(\out[1592]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1592]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_10 
       (.I0(padder_out_1[372]),
        .I1(out[308]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1356]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_11 
       (.I0(padder_out_1[512]),
        .I1(out[448]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1592]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_12 
       (.I0(padder_out_1[463]),
        .I1(out[399]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1527]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_13 
       (.I0(padder_out_1[256]),
        .I1(out[192]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1336]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1592]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[696] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1016] ),
        .I2(\f_permutation_l_/out_reg_n_0_[56] ),
        .I3(\f_permutation_l_/out_reg_n_0_[376] ),
        .O(\out[1592]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_2 
       (.I0(padder_out_1[180]),
        .I1(out[116]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1164]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1592]_i_3 
       (.I0(\out[1592]_i_6_n_0 ),
        .I1(padder_out_1[564]),
        .I2(out[500]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1592]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1419]),
        .O(\out[1592]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1592]_i_4 
       (.I0(\out[1550]_i_16_n_0 ),
        .I1(padder_out_1[501]),
        .I2(out[437]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1592]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1356]),
        .O(\out[1592]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1592]_i_5 
       (.I0(\f_permutation_l_/round_in [1592]),
        .I1(\f_permutation_l_/round_in [1527]),
        .I2(\out[1570]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[1592]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1592]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[908] ),
        .I1(padder_out_1[244]),
        .I2(out[180]),
        .I3(\f_permutation_l_/out_reg_n_0_[268] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[588] ),
        .O(\out[1592]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1592]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[779] ),
        .I1(padder_out_1[115]),
        .I2(out[51]),
        .I3(\f_permutation_l_/out_reg_n_0_[139] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[459] ),
        .O(\out[1592]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1592]_i_8 
       (.I0(padder_out_1[435]),
        .I1(out[371]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1419]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1592]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[716] ),
        .I1(padder_out_1[52]),
        .I2(\f_permutation_l_/out_reg_n_0_[1036] ),
        .I3(\f_permutation_l_/out_reg_n_0_[76] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[396] ),
        .O(\out[1592]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1593]_i_1 
       (.I0(\f_permutation_l_/round_in [1165]),
        .I1(\out[1593]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[782] ),
        .I3(\out[1593]_i_4_n_0 ),
        .I4(\out[1593]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1593]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_10 
       (.I0(padder_out_1[373]),
        .I1(out[309]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1357]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_11 
       (.I0(padder_out_1[513]),
        .I1(out[449]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1593]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_12 
       (.I0(padder_out_1[448]),
        .I1(out[384]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1528]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_13 
       (.I0(padder_out_1[257]),
        .I1(out[193]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1337]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1593]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[697] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1017] ),
        .I2(\f_permutation_l_/out_reg_n_0_[57] ),
        .I3(\f_permutation_l_/out_reg_n_0_[377] ),
        .O(\out[1593]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_2 
       (.I0(padder_out_1[181]),
        .I1(out[117]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1165]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1593]_i_3 
       (.I0(\out[1593]_i_6_n_0 ),
        .I1(padder_out_1[565]),
        .I2(out[501]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1593]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1420]),
        .O(\out[1593]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1593]_i_4 
       (.I0(\out[1551]_i_17_n_0 ),
        .I1(padder_out_1[502]),
        .I2(out[438]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1593]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1357]),
        .O(\out[1593]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1593]_i_5 
       (.I0(\f_permutation_l_/round_in [1593]),
        .I1(\f_permutation_l_/round_in [1528]),
        .I2(\out[1571]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[1593]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1593]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[909] ),
        .I1(padder_out_1[245]),
        .I2(out[181]),
        .I3(\f_permutation_l_/out_reg_n_0_[269] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[589] ),
        .O(\out[1593]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1593]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[780] ),
        .I1(padder_out_1[116]),
        .I2(out[52]),
        .I3(\f_permutation_l_/out_reg_n_0_[140] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[460] ),
        .O(\out[1593]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1593]_i_8 
       (.I0(padder_out_1[436]),
        .I1(out[372]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1420]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1593]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[717] ),
        .I1(padder_out_1[53]),
        .I2(\f_permutation_l_/out_reg_n_0_[1037] ),
        .I3(\f_permutation_l_/out_reg_n_0_[77] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[397] ),
        .O(\out[1593]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1594]_i_1 
       (.I0(\f_permutation_l_/round_in [1166]),
        .I1(\out[1594]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[783] ),
        .I3(\out[1594]_i_4_n_0 ),
        .I4(\out[1594]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1594]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_10 
       (.I0(padder_out_1[374]),
        .I1(out[310]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1358]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_11 
       (.I0(padder_out_1[514]),
        .I1(out[450]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1594]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_12 
       (.I0(padder_out_1[449]),
        .I1(out[385]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1529]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_13 
       (.I0(padder_out_1[258]),
        .I1(out[194]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1338]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1594]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[698] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1018] ),
        .I2(\f_permutation_l_/out_reg_n_0_[58] ),
        .I3(\f_permutation_l_/out_reg_n_0_[378] ),
        .O(\out[1594]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_2 
       (.I0(padder_out_1[182]),
        .I1(out[118]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1166]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1594]_i_3 
       (.I0(\out[1594]_i_6_n_0 ),
        .I1(padder_out_1[566]),
        .I2(out[502]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1594]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1421]),
        .O(\out[1594]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1594]_i_4 
       (.I0(\out[1552]_i_16_n_0 ),
        .I1(padder_out_1[503]),
        .I2(out[439]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1594]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1358]),
        .O(\out[1594]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1594]_i_5 
       (.I0(\f_permutation_l_/round_in [1594]),
        .I1(\f_permutation_l_/round_in [1529]),
        .I2(\out[1572]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[1594]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1594]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[910] ),
        .I1(padder_out_1[246]),
        .I2(out[182]),
        .I3(\f_permutation_l_/out_reg_n_0_[270] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[590] ),
        .O(\out[1594]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1594]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[781] ),
        .I1(padder_out_1[117]),
        .I2(out[53]),
        .I3(\f_permutation_l_/out_reg_n_0_[141] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[461] ),
        .O(\out[1594]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1594]_i_8 
       (.I0(padder_out_1[437]),
        .I1(out[373]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1421]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1594]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[718] ),
        .I1(padder_out_1[54]),
        .I2(\f_permutation_l_/out_reg_n_0_[1038] ),
        .I3(\f_permutation_l_/out_reg_n_0_[78] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[398] ),
        .O(\out[1594]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1595]_i_1 
       (.I0(\f_permutation_l_/round_in [1167]),
        .I1(\out[1595]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[784] ),
        .I3(\out[1595]_i_4_n_0 ),
        .I4(\out[1595]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1595]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_10 
       (.I0(padder_out_1[375]),
        .I1(out[311]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1359]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_11 
       (.I0(padder_out_1[515]),
        .I1(out[451]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1595]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_12 
       (.I0(padder_out_1[450]),
        .I1(out[386]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1530]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_13 
       (.I0(padder_out_1[259]),
        .I1(out[195]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1339]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1595]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[699] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1019] ),
        .I2(\f_permutation_l_/out_reg_n_0_[59] ),
        .I3(\f_permutation_l_/out_reg_n_0_[379] ),
        .O(\out[1595]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_2 
       (.I0(padder_out_1[183]),
        .I1(out[119]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1167]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1595]_i_3 
       (.I0(\out[1595]_i_6_n_0 ),
        .I1(padder_out_1[567]),
        .I2(out[503]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1595]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1422]),
        .O(\out[1595]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1595]_i_4 
       (.I0(\out[1553]_i_16_n_0 ),
        .I1(padder_out_1[488]),
        .I2(out[424]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1595]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1359]),
        .O(\out[1595]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1595]_i_5 
       (.I0(\f_permutation_l_/round_in [1595]),
        .I1(\f_permutation_l_/round_in [1530]),
        .I2(\out[1573]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[1595]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1595]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[911] ),
        .I1(padder_out_1[247]),
        .I2(out[183]),
        .I3(\f_permutation_l_/out_reg_n_0_[271] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[591] ),
        .O(\out[1595]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1595]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[782] ),
        .I1(padder_out_1[118]),
        .I2(out[54]),
        .I3(\f_permutation_l_/out_reg_n_0_[142] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[462] ),
        .O(\out[1595]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1595]_i_8 
       (.I0(padder_out_1[438]),
        .I1(out[374]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1422]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1595]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[719] ),
        .I1(padder_out_1[55]),
        .I2(\f_permutation_l_/out_reg_n_0_[1039] ),
        .I3(\f_permutation_l_/out_reg_n_0_[79] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[399] ),
        .O(\out[1595]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1596]_i_1 
       (.I0(\f_permutation_l_/round_in [1168]),
        .I1(\out[1596]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[785] ),
        .I3(\out[1596]_i_4_n_0 ),
        .I4(\out[1596]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1596]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_10 
       (.I0(padder_out_1[360]),
        .I1(out[296]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1360]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_11 
       (.I0(padder_out_1[516]),
        .I1(out[452]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1596]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_12 
       (.I0(padder_out_1[451]),
        .I1(out[387]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1531]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_13 
       (.I0(padder_out_1[260]),
        .I1(out[196]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1340]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1596]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[700] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1020] ),
        .I2(\f_permutation_l_/out_reg_n_0_[60] ),
        .I3(\f_permutation_l_/out_reg_n_0_[380] ),
        .O(\out[1596]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_2 
       (.I0(padder_out_1[168]),
        .I1(out[104]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1168]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1596]_i_3 
       (.I0(\out[1596]_i_6_n_0 ),
        .I1(padder_out_1[552]),
        .I2(out[488]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1596]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1423]),
        .O(\out[1596]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1596]_i_4 
       (.I0(\out[1554]_i_16_n_0 ),
        .I1(padder_out_1[489]),
        .I2(out[425]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1596]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1360]),
        .O(\out[1596]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1596]_i_5 
       (.I0(\f_permutation_l_/round_in [1596]),
        .I1(\f_permutation_l_/round_in [1531]),
        .I2(\out[1574]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[1596]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1596]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[912] ),
        .I1(padder_out_1[232]),
        .I2(out[168]),
        .I3(\f_permutation_l_/out_reg_n_0_[272] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[592] ),
        .O(\out[1596]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1596]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[783] ),
        .I1(padder_out_1[119]),
        .I2(out[55]),
        .I3(\f_permutation_l_/out_reg_n_0_[143] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[463] ),
        .O(\out[1596]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1596]_i_8 
       (.I0(padder_out_1[439]),
        .I1(out[375]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1423]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1596]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[720] ),
        .I1(padder_out_1[40]),
        .I2(\f_permutation_l_/out_reg_n_0_[1040] ),
        .I3(\f_permutation_l_/out_reg_n_0_[80] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[400] ),
        .O(\out[1596]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1597]_i_1 
       (.I0(\f_permutation_l_/round_in [1169]),
        .I1(\out[1597]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[786] ),
        .I3(\out[1597]_i_4_n_0 ),
        .I4(\out[1597]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1597]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_10 
       (.I0(padder_out_1[361]),
        .I1(out[297]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1361]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_11 
       (.I0(padder_out_1[517]),
        .I1(out[453]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1597]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_12 
       (.I0(padder_out_1[452]),
        .I1(out[388]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1532]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_13 
       (.I0(padder_out_1[261]),
        .I1(out[197]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1341]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1597]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[701] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1021] ),
        .I2(\f_permutation_l_/out_reg_n_0_[61] ),
        .I3(\f_permutation_l_/out_reg_n_0_[381] ),
        .O(\out[1597]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_2 
       (.I0(padder_out_1[169]),
        .I1(out[105]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1169]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1597]_i_3 
       (.I0(\out[1597]_i_6_n_0 ),
        .I1(padder_out_1[553]),
        .I2(out[489]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1597]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1424]),
        .O(\out[1597]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1597]_i_4 
       (.I0(\out[1555]_i_16_n_0 ),
        .I1(padder_out_1[490]),
        .I2(out[426]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1597]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1361]),
        .O(\out[1597]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1597]_i_5 
       (.I0(\f_permutation_l_/round_in [1597]),
        .I1(\f_permutation_l_/round_in [1532]),
        .I2(\out[1575]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[1597]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1597]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[913] ),
        .I1(padder_out_1[233]),
        .I2(out[169]),
        .I3(\f_permutation_l_/out_reg_n_0_[273] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[593] ),
        .O(\out[1597]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1597]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[784] ),
        .I1(padder_out_1[104]),
        .I2(out[40]),
        .I3(\f_permutation_l_/out_reg_n_0_[144] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[464] ),
        .O(\out[1597]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1597]_i_8 
       (.I0(padder_out_1[424]),
        .I1(out[360]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1424]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1597]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[721] ),
        .I1(padder_out_1[41]),
        .I2(\f_permutation_l_/out_reg_n_0_[1041] ),
        .I3(\f_permutation_l_/out_reg_n_0_[81] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[401] ),
        .O(\out[1597]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[1598]_i_1 
       (.I0(\f_permutation_l_/round_in [1170]),
        .I1(\out[1598]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[787] ),
        .I3(\out[1598]_i_4_n_0 ),
        .I4(\out[1598]_i_5_n_0 ),
        .O(\f_permutation_l_/round_out [1598]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_10 
       (.I0(padder_out_1[362]),
        .I1(out[298]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1362]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_11 
       (.I0(padder_out_1[518]),
        .I1(out[454]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1598]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_12 
       (.I0(padder_out_1[453]),
        .I1(out[389]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1533]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_13 
       (.I0(padder_out_1[262]),
        .I1(out[198]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1342]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1598]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[702] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1022] ),
        .I2(\f_permutation_l_/out_reg_n_0_[62] ),
        .I3(\f_permutation_l_/out_reg_n_0_[382] ),
        .O(\out[1598]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_2 
       (.I0(padder_out_1[170]),
        .I1(out[106]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1170]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h69A5965A965A69A5)) 
    \out[1598]_i_3 
       (.I0(\out[1598]_i_6_n_0 ),
        .I1(padder_out_1[554]),
        .I2(out[490]),
        .I3(\out[1542]_i_8_n_0 ),
        .I4(\out[1598]_i_7_n_0 ),
        .I5(\f_permutation_l_/round_in [1425]),
        .O(\out[1598]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1598]_i_4 
       (.I0(\out[1556]_i_16_n_0 ),
        .I1(padder_out_1[491]),
        .I2(out[427]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1598]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1362]),
        .O(\out[1598]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1598]_i_5 
       (.I0(\f_permutation_l_/round_in [1598]),
        .I1(\f_permutation_l_/round_in [1533]),
        .I2(\out[1576]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[1598]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1598]_i_6 
       (.I0(\f_permutation_l_/out_reg_n_0_[914] ),
        .I1(padder_out_1[234]),
        .I2(out[170]),
        .I3(\f_permutation_l_/out_reg_n_0_[274] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[594] ),
        .O(\out[1598]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1598]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[785] ),
        .I1(padder_out_1[105]),
        .I2(out[41]),
        .I3(\f_permutation_l_/out_reg_n_0_[145] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[465] ),
        .O(\out[1598]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1598]_i_8 
       (.I0(padder_out_1[425]),
        .I1(out[361]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1425]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1598]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[722] ),
        .I1(padder_out_1[42]),
        .I2(\f_permutation_l_/out_reg_n_0_[1042] ),
        .I3(\f_permutation_l_/out_reg_n_0_[82] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[402] ),
        .O(\out[1598]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h14EBEB14)) 
    \out[1599]_i_1 
       (.I0(\out[1599]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[788] ),
        .I2(\out[1599]_i_3_n_0 ),
        .I3(\out[1599]_i_4_n_0 ),
        .I4(\f_permutation_l_/rc [63]),
        .O(\f_permutation_l_/round_out [1599]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1599]_i_10 
       (.I0(padder_out_1[363]),
        .I1(out[299]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1363]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1599]_i_11 
       (.I0(padder_out_1[519]),
        .I1(out[455]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1599]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1599]_i_12 
       (.I0(padder_out_1[454]),
        .I1(out[390]),
        .I2(\out[1415]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1534]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1599]_i_13 
       (.I0(padder_out_1[263]),
        .I1(out[199]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1343]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h6996)) 
    \out[1599]_i_14 
       (.I0(\f_permutation_l_/out_reg_n_0_[703] ),
        .I1(\f_permutation_l_/out_reg_n_0_[1023] ),
        .I2(\f_permutation_l_/out_reg_n_0_[63] ),
        .I3(\f_permutation_l_/out_reg_n_0_[383] ),
        .O(\out[1599]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1599]_i_15 
       (.I0(\out[1543]_i_21_n_0 ),
        .I1(\f_permutation_l_/i_reg_n_0_[1] ),
        .I2(\f_permutation_l_/i_reg_n_0_[12] ),
        .I3(\f_permutation_l_/i_reg_n_0_[14] ),
        .I4(\f_permutation_l_/i_reg_n_0_[15] ),
        .I5(\f_permutation_l_/i_reg_n_0_[16] ),
        .O(\out[1599]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1599]_i_2 
       (.I0(\f_permutation_l_/round_in [1171]),
        .I1(\f_permutation_l_/round_in [1426]),
        .I2(\out[1599]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1555]),
        .I4(\out[1599]_i_8_n_0 ),
        .O(\out[1599]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h965A69A569A5965A)) 
    \out[1599]_i_3 
       (.I0(\out[1557]_i_15_n_0 ),
        .I1(padder_out_1[492]),
        .I2(out[428]),
        .I3(\out[1543]_i_12_n_0 ),
        .I4(\out[1599]_i_9_n_0 ),
        .I5(\f_permutation_l_/round_in [1363]),
        .O(\out[1599]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[1599]_i_4 
       (.I0(\f_permutation_l_/round_in [1599]),
        .I1(\f_permutation_l_/round_in [1534]),
        .I2(\out[1577]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[1599]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \out[1599]_i_5 
       (.I0(\out[1599]_i_15_n_0 ),
        .I1(\f_permutation_l_/i_reg_n_0_[18] ),
        .I2(\f_permutation_l_/i_reg_n_0_[13] ),
        .I3(\f_permutation_l_/i_reg_n_0_[6] ),
        .I4(\f_permutation_l_/i_reg_n_0_[2] ),
        .I5(\f_permutation_l_/p_0_in ),
        .O(\f_permutation_l_/rc [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[1599]_i_6 
       (.I0(padder_out_1[426]),
        .I1(out[362]),
        .I2(\out[1556]_i_7_n_0 ),
        .O(\f_permutation_l_/round_in [1426]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1599]_i_7 
       (.I0(\f_permutation_l_/out_reg_n_0_[786] ),
        .I1(padder_out_1[106]),
        .I2(out[42]),
        .I3(\f_permutation_l_/out_reg_n_0_[146] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[466] ),
        .O(\out[1599]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1599]_i_8 
       (.I0(\f_permutation_l_/out_reg_n_0_[915] ),
        .I1(padder_out_1[235]),
        .I2(out[171]),
        .I3(\f_permutation_l_/out_reg_n_0_[275] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[595] ),
        .O(\out[1599]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h96695AA56996A55A)) 
    \out[1599]_i_9 
       (.I0(\f_permutation_l_/out_reg_n_0_[723] ),
        .I1(padder_out_1[43]),
        .I2(\f_permutation_l_/out_reg_n_0_[1043] ),
        .I3(\f_permutation_l_/out_reg_n_0_[83] ),
        .I4(update__0_i_1_n_0),
        .I5(\f_permutation_l_/out_reg_n_0_[403] ),
        .O(\out[1599]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[159]_i_1 
       (.I0(\out[1414]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[696] ),
        .I2(\out[159]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[221] ),
        .I4(\out[1545]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [159]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[159]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[630] ),
        .I1(\f_permutation_l_/round_in [1525]),
        .I2(\out[1568]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[159]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[15]_i_1 
       (.I0(\out[1593]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[205] ),
        .I2(\out[271]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1048]),
        .I4(\out[1517]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[160]_i_1 
       (.I0(\out[1415]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[697] ),
        .I2(\out[160]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[222] ),
        .I4(\out[1546]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [160]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[160]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[631] ),
        .I1(\f_permutation_l_/round_in [1526]),
        .I2(\out[1569]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[160]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[161]_i_1 
       (.I0(\out[1416]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[698] ),
        .I2(\out[161]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[223] ),
        .I4(\out[1547]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [161]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[161]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[632] ),
        .I1(\f_permutation_l_/round_in [1527]),
        .I2(\out[1570]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[161]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[162]_i_1 
       (.I0(\out[1417]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[699] ),
        .I2(\out[162]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[224] ),
        .I4(\out[1548]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [162]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[162]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[633] ),
        .I1(\f_permutation_l_/round_in [1528]),
        .I2(\out[1571]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[162]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[163]_i_1 
       (.I0(\out[1418]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[700] ),
        .I2(\out[163]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[225] ),
        .I4(\out[1549]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [163]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[163]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[634] ),
        .I1(\f_permutation_l_/round_in [1529]),
        .I2(\out[1572]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[163]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[164]_i_1 
       (.I0(\out[1419]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[701] ),
        .I2(\out[164]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[226] ),
        .I4(\out[1550]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [164]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[164]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[635] ),
        .I1(\f_permutation_l_/round_in [1530]),
        .I2(\out[1573]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[164]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[165]_i_1 
       (.I0(\out[1420]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[702] ),
        .I2(\out[165]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[227] ),
        .I4(\out[1295]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [165]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[165]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[636] ),
        .I1(\f_permutation_l_/round_in [1531]),
        .I2(\out[1574]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[165]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[166]_i_1 
       (.I0(\out[1421]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[703] ),
        .I2(\out[166]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[228] ),
        .I4(\out[1552]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [166]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[166]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[637] ),
        .I1(\f_permutation_l_/round_in [1532]),
        .I2(\out[1575]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[166]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[167]_i_1 
       (.I0(\out[1422]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[640] ),
        .I2(\out[167]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[229] ),
        .I4(\out[1553]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [167]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[167]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[638] ),
        .I1(\f_permutation_l_/round_in [1533]),
        .I2(\out[1576]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[167]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[168]_i_1 
       (.I0(\out[1423]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[641] ),
        .I2(\out[168]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[230] ),
        .I4(\out[1554]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [168]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[168]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[639] ),
        .I1(\f_permutation_l_/round_in [1534]),
        .I2(\out[1577]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[168]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[169]_i_1 
       (.I0(\out[1424]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[642] ),
        .I2(\out[169]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[231] ),
        .I4(\out[1555]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [169]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[169]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[576] ),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[169]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[16]_i_1 
       (.I0(\out[1594]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[206] ),
        .I2(\out[272]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1049]),
        .I4(\out[1518]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[170]_i_1 
       (.I0(\out[1425]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[643] ),
        .I2(\out[170]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[232] ),
        .I4(\out[1556]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [170]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[170]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[577] ),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[170]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[171]_i_1 
       (.I0(\out[1426]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[644] ),
        .I2(\out[171]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[233] ),
        .I4(\out[1557]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [171]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[171]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[578] ),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[171]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[172]_i_1 
       (.I0(\out[1427]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[645] ),
        .I2(\out[172]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[234] ),
        .I4(\out[1558]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [172]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[172]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[579] ),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[172]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[173]_i_1 
       (.I0(\out[1428]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[646] ),
        .I2(\out[173]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[235] ),
        .I4(\out[1559]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [173]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[173]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[580] ),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[173]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[174]_i_1 
       (.I0(\out[1429]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[647] ),
        .I2(\out[174]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[236] ),
        .I4(\out[1560]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [174]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[174]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[581] ),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[174]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[175]_i_1 
       (.I0(\out[1430]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[648] ),
        .I2(\out[175]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[237] ),
        .I4(\out[1561]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [175]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[175]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[582] ),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[175]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[176]_i_1 
       (.I0(\out[1431]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[649] ),
        .I2(\out[176]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[238] ),
        .I4(\out[1562]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [176]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[176]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[583] ),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[176]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[177]_i_1 
       (.I0(\out[1432]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[650] ),
        .I2(\out[177]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[239] ),
        .I4(\out[1563]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [177]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[177]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[584] ),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[177]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[178]_i_1 
       (.I0(\out[1433]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[651] ),
        .I2(\out[178]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[240] ),
        .I4(\out[1564]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [178]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[178]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[585] ),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[178]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[179]_i_1 
       (.I0(\out[1434]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[652] ),
        .I2(\out[179]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[241] ),
        .I4(\out[1565]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [179]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[179]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[586] ),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[179]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[17]_i_1 
       (.I0(\out[1595]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[207] ),
        .I2(\out[273]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1050]),
        .I4(\out[1519]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[180]_i_1 
       (.I0(\out[1435]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[653] ),
        .I2(\out[180]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[242] ),
        .I4(\out[1566]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [180]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[180]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[587] ),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[180]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[181]_i_1 
       (.I0(\out[1436]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[654] ),
        .I2(\out[181]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[243] ),
        .I4(\out[1311]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [181]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[181]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[588] ),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[181]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[182]_i_1 
       (.I0(\out[1437]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[655] ),
        .I2(\out[182]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[244] ),
        .I4(\out[1568]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [182]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[182]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[589] ),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[182]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[183]_i_1 
       (.I0(\out[1438]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[656] ),
        .I2(\out[183]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[245] ),
        .I4(\out[1569]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [183]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[183]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[590] ),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[183]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[184]_i_1 
       (.I0(\out[1439]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[657] ),
        .I2(\out[184]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[246] ),
        .I4(\out[1570]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [184]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[184]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[591] ),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[184]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[185]_i_1 
       (.I0(\out[1440]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[658] ),
        .I2(\out[185]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[247] ),
        .I4(\out[1571]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [185]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[185]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[592] ),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[185]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[186]_i_1 
       (.I0(\out[1441]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[659] ),
        .I2(\out[186]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[248] ),
        .I4(\out[1572]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [186]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[186]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[593] ),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[186]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[187]_i_1 
       (.I0(\out[1442]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[660] ),
        .I2(\out[187]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[249] ),
        .I4(\out[1573]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [187]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[187]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[594] ),
        .I1(\f_permutation_l_/round_in [1298]),
        .I2(\out[1554]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[187]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[188]_i_1 
       (.I0(\out[1443]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[661] ),
        .I2(\out[188]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[250] ),
        .I4(\out[1574]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [188]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[188]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[595] ),
        .I1(\f_permutation_l_/round_in [1299]),
        .I2(\out[1555]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[188]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[189]_i_1 
       (.I0(\out[1444]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[662] ),
        .I2(\out[189]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[251] ),
        .I4(\out[1575]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [189]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[189]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[596] ),
        .I1(\f_permutation_l_/round_in [1300]),
        .I2(\out[1556]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[189]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[18]_i_1 
       (.I0(\out[1596]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[208] ),
        .I2(\out[274]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1051]),
        .I4(\out[1520]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[190]_i_1 
       (.I0(\out[1445]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[663] ),
        .I2(\out[190]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[252] ),
        .I4(\out[1576]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [190]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[190]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[597] ),
        .I1(\f_permutation_l_/round_in [1301]),
        .I2(\out[1557]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[190]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[191]_i_1 
       (.I0(\out[1446]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[664] ),
        .I2(\out[191]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[253] ),
        .I4(\out[1577]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [191]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[191]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[598] ),
        .I1(\out[1536]_i_14_n_0 ),
        .I2(\f_permutation_l_/round_in [1493]),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[191]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[192]_i_1 
       (.I0(\out[192]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[665] ),
        .I2(\out[1447]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[599] ),
        .I4(\out[1242]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [192]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[192]_i_2 
       (.I0(\f_permutation_l_/round_in [1033]),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1417]),
        .I4(\out[1590]_i_7_n_0 ),
        .O(\out[192]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[193]_i_1 
       (.I0(\out[193]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[666] ),
        .I2(\out[1448]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[600] ),
        .I4(\out[1243]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [193]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[193]_i_2 
       (.I0(\f_permutation_l_/round_in [1034]),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1418]),
        .I4(\out[1591]_i_7_n_0 ),
        .O(\out[193]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[194]_i_1 
       (.I0(\out[194]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[667] ),
        .I2(\out[1449]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[601] ),
        .I4(\out[1244]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [194]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[194]_i_2 
       (.I0(\f_permutation_l_/round_in [1035]),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1419]),
        .I4(\out[1592]_i_7_n_0 ),
        .O(\out[194]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[195]_i_1 
       (.I0(\out[195]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[668] ),
        .I2(\out[1450]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[602] ),
        .I4(\out[1245]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [195]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[195]_i_2 
       (.I0(\f_permutation_l_/round_in [1036]),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1420]),
        .I4(\out[1593]_i_7_n_0 ),
        .O(\out[195]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[196]_i_1 
       (.I0(\out[196]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[669] ),
        .I2(\out[1451]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[603] ),
        .I4(\out[1246]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [196]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[196]_i_2 
       (.I0(\f_permutation_l_/round_in [1037]),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1421]),
        .I4(\out[1594]_i_7_n_0 ),
        .O(\out[196]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[197]_i_1 
       (.I0(\out[197]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[670] ),
        .I2(\out[1452]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[604] ),
        .I4(\out[1247]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [197]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[197]_i_2 
       (.I0(\f_permutation_l_/round_in [1038]),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1422]),
        .I4(\out[1595]_i_7_n_0 ),
        .O(\out[197]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[198]_i_1 
       (.I0(\out[198]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[671] ),
        .I2(\out[1453]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[605] ),
        .I4(\out[1248]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [198]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[198]_i_2 
       (.I0(\f_permutation_l_/round_in [1039]),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1423]),
        .I4(\out[1596]_i_7_n_0 ),
        .O(\out[198]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[199]_i_1 
       (.I0(\out[199]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[672] ),
        .I2(\out[1454]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[606] ),
        .I4(\out[1249]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [199]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[199]_i_2 
       (.I0(\f_permutation_l_/round_in [1040]),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1424]),
        .I4(\out[1597]_i_7_n_0 ),
        .O(\out[199]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[19]_i_1 
       (.I0(\out[1597]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[209] ),
        .I2(\out[275]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1052]),
        .I4(\out[1521]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[1]_i_1 
       (.I0(\out[1579]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[255] ),
        .I2(\out[257]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1034]),
        .I4(\out[1503]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[200]_i_1 
       (.I0(\out[200]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[673] ),
        .I2(\out[1455]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[607] ),
        .I4(\out[1250]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [200]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[200]_i_2 
       (.I0(\f_permutation_l_/round_in [1041]),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1425]),
        .I4(\out[1598]_i_7_n_0 ),
        .O(\out[200]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[201]_i_1 
       (.I0(\out[201]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[674] ),
        .I2(\out[1456]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[608] ),
        .I4(\out[1251]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [201]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[201]_i_2 
       (.I0(\f_permutation_l_/round_in [1042]),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\out[1599]_i_7_n_0 ),
        .I4(\f_permutation_l_/round_in [1426]),
        .O(\out[201]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[202]_i_1 
       (.I0(\out[202]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[675] ),
        .I2(\out[1457]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[609] ),
        .I4(\out[1252]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [202]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[202]_i_2 
       (.I0(\f_permutation_l_/round_in [1043]),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\out[1554]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1298]),
        .O(\out[202]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[203]_i_1 
       (.I0(\out[203]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[676] ),
        .I2(\out[1458]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[610] ),
        .I4(\out[1253]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [203]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[203]_i_2 
       (.I0(\f_permutation_l_/round_in [1044]),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\out[1555]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1299]),
        .O(\out[203]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[204]_i_1 
       (.I0(\out[204]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[677] ),
        .I2(\out[1459]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[611] ),
        .I4(\out[1254]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [204]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[204]_i_2 
       (.I0(\f_permutation_l_/round_in [1045]),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\out[1556]_i_14_n_0 ),
        .I4(\f_permutation_l_/round_in [1300]),
        .O(\out[204]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[205]_i_1 
       (.I0(\out[205]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[678] ),
        .I2(\out[1460]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[612] ),
        .I4(\out[1255]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [205]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[205]_i_2 
       (.I0(\f_permutation_l_/round_in [1046]),
        .I1(\f_permutation_l_/round_in [1430]),
        .I2(\out[1539]_i_9_n_0 ),
        .I3(\out[1557]_i_13_n_0 ),
        .I4(\f_permutation_l_/round_in [1301]),
        .O(\out[205]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[206]_i_1 
       (.I0(\out[206]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[679] ),
        .I2(\out[1461]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[613] ),
        .I4(\out[1256]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [206]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[206]_i_2 
       (.I0(\f_permutation_l_/round_in [1047]),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[206]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[207]_i_1 
       (.I0(\out[207]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[680] ),
        .I2(\out[1462]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[614] ),
        .I4(\out[1257]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [207]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[207]_i_2 
       (.I0(\f_permutation_l_/round_in [1048]),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[207]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[208]_i_1 
       (.I0(\out[208]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[681] ),
        .I2(\out[1463]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[615] ),
        .I4(\out[1258]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [208]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[208]_i_2 
       (.I0(\f_permutation_l_/round_in [1049]),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[208]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[209]_i_1 
       (.I0(\out[209]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[682] ),
        .I2(\out[1464]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[616] ),
        .I4(\out[1259]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [209]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[209]_i_2 
       (.I0(\f_permutation_l_/round_in [1050]),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[209]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[20]_i_1 
       (.I0(\out[1598]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[210] ),
        .I2(\out[276]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1053]),
        .I4(\out[1522]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[210]_i_1 
       (.I0(\out[210]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[683] ),
        .I2(\out[1465]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[617] ),
        .I4(\out[1260]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [210]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[210]_i_2 
       (.I0(\f_permutation_l_/round_in [1051]),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[210]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[211]_i_1 
       (.I0(\out[211]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[684] ),
        .I2(\out[1466]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[618] ),
        .I4(\out[1261]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [211]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[211]_i_2 
       (.I0(\f_permutation_l_/round_in [1052]),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[211]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[212]_i_1 
       (.I0(\out[212]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[685] ),
        .I2(\out[1467]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[619] ),
        .I4(\out[1262]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [212]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[212]_i_2 
       (.I0(\f_permutation_l_/round_in [1053]),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[212]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[213]_i_1 
       (.I0(\out[213]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[686] ),
        .I2(\out[1468]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[620] ),
        .I4(\out[1263]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [213]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[213]_i_2 
       (.I0(\f_permutation_l_/round_in [1054]),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[213]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[214]_i_1 
       (.I0(\out[214]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[687] ),
        .I2(\out[1469]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[621] ),
        .I4(\out[1264]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [214]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[214]_i_2 
       (.I0(\f_permutation_l_/round_in [1055]),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[214]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[215]_i_1 
       (.I0(\out[215]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[688] ),
        .I2(\out[1470]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[622] ),
        .I4(\out[1265]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [215]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[215]_i_2 
       (.I0(\f_permutation_l_/round_in [1056]),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[215]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[216]_i_1 
       (.I0(\out[216]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[689] ),
        .I2(\out[1471]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[623] ),
        .I4(\out[1266]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [216]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[216]_i_2 
       (.I0(\f_permutation_l_/round_in [1057]),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[216]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[217]_i_1 
       (.I0(\out[217]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[690] ),
        .I2(\out[1408]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[624] ),
        .I4(\out[1267]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [217]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[217]_i_2 
       (.I0(\f_permutation_l_/round_in [1058]),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[217]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[218]_i_1 
       (.I0(\out[218]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[691] ),
        .I2(\out[1409]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[625] ),
        .I4(\out[1268]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [218]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[218]_i_2 
       (.I0(\f_permutation_l_/round_in [1059]),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[218]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[219]_i_1 
       (.I0(\out[219]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[692] ),
        .I2(\out[1410]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[626] ),
        .I4(\out[1269]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [219]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[219]_i_2 
       (.I0(\f_permutation_l_/round_in [1060]),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[219]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[21]_i_1 
       (.I0(\out[1343]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[211] ),
        .I2(\out[277]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1054]),
        .I4(\out[1523]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[220]_i_1 
       (.I0(\out[220]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[693] ),
        .I2(\out[1411]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[627] ),
        .I4(\out[1270]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [220]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[220]_i_2 
       (.I0(\f_permutation_l_/round_in [1061]),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[220]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[221]_i_1 
       (.I0(\out[221]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[694] ),
        .I2(\out[1412]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[628] ),
        .I4(\out[1271]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [221]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[221]_i_2 
       (.I0(\f_permutation_l_/round_in [1062]),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[221]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[222]_i_1 
       (.I0(\out[222]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[695] ),
        .I2(\out[1413]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[629] ),
        .I4(\out[1272]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [222]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[222]_i_2 
       (.I0(\f_permutation_l_/round_in [1063]),
        .I1(\f_permutation_l_/round_in [1447]),
        .I2(\out[1556]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[222]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[223]_i_1 
       (.I0(\out[223]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[696] ),
        .I2(\out[1414]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[630] ),
        .I4(\out[1273]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [223]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[223]_i_2 
       (.I0(\f_permutation_l_/round_in [1064]),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[223]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[224]_i_1 
       (.I0(\out[224]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[697] ),
        .I2(\out[1415]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[631] ),
        .I4(\out[1274]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [224]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[224]_i_2 
       (.I0(\f_permutation_l_/round_in [1065]),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[224]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[225]_i_1 
       (.I0(\out[225]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[698] ),
        .I2(\out[1416]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[632] ),
        .I4(\out[1275]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [225]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[225]_i_2 
       (.I0(\f_permutation_l_/round_in [1066]),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[225]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[226]_i_1 
       (.I0(\out[226]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[699] ),
        .I2(\out[1417]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[633] ),
        .I4(\out[1276]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [226]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[226]_i_2 
       (.I0(\f_permutation_l_/round_in [1067]),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[226]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[227]_i_1 
       (.I0(\out[227]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[700] ),
        .I2(\out[1418]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[634] ),
        .I4(\out[1277]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [227]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[227]_i_2 
       (.I0(\f_permutation_l_/round_in [1068]),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[227]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[228]_i_1 
       (.I0(\out[228]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[701] ),
        .I2(\out[1419]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[635] ),
        .I4(\out[1278]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [228]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[228]_i_2 
       (.I0(\f_permutation_l_/round_in [1069]),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[228]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[229]_i_1 
       (.I0(\out[229]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[702] ),
        .I2(\out[1420]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[636] ),
        .I4(\out[1279]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [229]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[229]_i_2 
       (.I0(\f_permutation_l_/round_in [1070]),
        .I1(\f_permutation_l_/round_in [1454]),
        .I2(\out[1563]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[229]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[22]_i_1 
       (.I0(\out[1280]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[212] ),
        .I2(\out[278]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1055]),
        .I4(\out[1524]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[230]_i_1 
       (.I0(\out[230]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[703] ),
        .I2(\out[1421]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[637] ),
        .I4(\out[1216]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [230]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[230]_i_2 
       (.I0(\f_permutation_l_/round_in [1071]),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[230]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[231]_i_1 
       (.I0(\out[231]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[640] ),
        .I2(\out[1422]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[638] ),
        .I4(\out[1217]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [231]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[231]_i_2 
       (.I0(\f_permutation_l_/round_in [1072]),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[231]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[232]_i_1 
       (.I0(\out[232]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[641] ),
        .I2(\out[1423]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[639] ),
        .I4(\out[1218]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [232]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[232]_i_2 
       (.I0(\f_permutation_l_/round_in [1073]),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[232]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[233]_i_1 
       (.I0(\out[233]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[642] ),
        .I2(\out[1424]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[576] ),
        .I4(\out[1219]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [233]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[233]_i_2 
       (.I0(\f_permutation_l_/round_in [1074]),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[233]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[234]_i_1 
       (.I0(\out[234]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[643] ),
        .I2(\out[1425]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[577] ),
        .I4(\out[1220]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [234]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[234]_i_2 
       (.I0(\f_permutation_l_/round_in [1075]),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[234]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[235]_i_1 
       (.I0(\out[235]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[644] ),
        .I2(\out[1426]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[578] ),
        .I4(\out[1221]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [235]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[235]_i_2 
       (.I0(\f_permutation_l_/round_in [1076]),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[235]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[236]_i_1 
       (.I0(\out[236]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[645] ),
        .I2(\out[1427]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[579] ),
        .I4(\out[1539]_i_6_n_0 ),
        .O(\f_permutation_l_/round_out [236]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[236]_i_2 
       (.I0(\f_permutation_l_/round_in [1077]),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[236]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[237]_i_1 
       (.I0(\out[237]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[646] ),
        .I2(\out[1428]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[580] ),
        .I4(\out[1223]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [237]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[237]_i_2 
       (.I0(\f_permutation_l_/round_in [1078]),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[237]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[238]_i_1 
       (.I0(\out[238]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[647] ),
        .I2(\out[1429]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[581] ),
        .I4(\out[1224]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [238]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[238]_i_2 
       (.I0(\f_permutation_l_/round_in [1079]),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[238]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[239]_i_1 
       (.I0(\out[239]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[648] ),
        .I2(\out[1430]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[582] ),
        .I4(\out[1225]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [239]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[239]_i_2 
       (.I0(\f_permutation_l_/round_in [1080]),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[239]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[23]_i_1 
       (.I0(\out[1281]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[213] ),
        .I2(\out[279]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1056]),
        .I4(\out[1525]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[240]_i_1 
       (.I0(\out[240]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[649] ),
        .I2(\out[1431]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[583] ),
        .I4(\out[1226]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [240]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[240]_i_2 
       (.I0(\f_permutation_l_/round_in [1081]),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[240]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[241]_i_1 
       (.I0(\out[241]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[650] ),
        .I2(\out[1432]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[584] ),
        .I4(\out[1227]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [241]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[241]_i_2 
       (.I0(\f_permutation_l_/round_in [1082]),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[241]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[242]_i_1 
       (.I0(\out[242]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[651] ),
        .I2(\out[1433]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[585] ),
        .I4(\out[1228]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [242]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[242]_i_2 
       (.I0(\f_permutation_l_/round_in [1083]),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[242]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[243]_i_1 
       (.I0(\out[243]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[652] ),
        .I2(\out[1434]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[586] ),
        .I4(\out[1229]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [243]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[243]_i_2 
       (.I0(\f_permutation_l_/round_in [1084]),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[243]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[244]_i_1 
       (.I0(\out[244]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[653] ),
        .I2(\out[1435]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[587] ),
        .I4(\out[1230]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [244]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[244]_i_2 
       (.I0(\f_permutation_l_/round_in [1085]),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[244]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[245]_i_1 
       (.I0(\out[245]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[654] ),
        .I2(\out[1436]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[588] ),
        .I4(\out[1231]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [245]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[245]_i_2 
       (.I0(\f_permutation_l_/round_in [1086]),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[245]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[246]_i_1 
       (.I0(\out[246]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[655] ),
        .I2(\out[1437]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[589] ),
        .I4(\out[1232]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [246]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[246]_i_2 
       (.I0(\f_permutation_l_/round_in [1087]),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[246]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[247]_i_1 
       (.I0(\out[247]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[656] ),
        .I2(\out[1438]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[590] ),
        .I4(\out[1233]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [247]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[247]_i_2 
       (.I0(\f_permutation_l_/round_in [1024]),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[247]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[248]_i_1 
       (.I0(\out[248]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[657] ),
        .I2(\out[1439]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[591] ),
        .I4(\out[1234]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [248]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[248]_i_2 
       (.I0(\f_permutation_l_/round_in [1025]),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1409]),
        .I4(\out[1582]_i_7_n_0 ),
        .O(\out[248]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[249]_i_1 
       (.I0(\out[249]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[658] ),
        .I2(\out[1440]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[592] ),
        .I4(\out[1235]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [249]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[249]_i_2 
       (.I0(\f_permutation_l_/round_in [1026]),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1410]),
        .I4(\out[1583]_i_7_n_0 ),
        .O(\out[249]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[24]_i_1 
       (.I0(\out[1538]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[214] ),
        .I2(\out[280]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1057]),
        .I4(\out[1526]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[250]_i_1 
       (.I0(\out[250]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[659] ),
        .I2(\out[1441]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[593] ),
        .I4(\out[1236]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [250]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[250]_i_2 
       (.I0(\f_permutation_l_/round_in [1027]),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1411]),
        .I4(\out[1584]_i_7_n_0 ),
        .O(\out[250]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[251]_i_1 
       (.I0(\out[251]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[660] ),
        .I2(\out[1442]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[594] ),
        .I4(\out[1237]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [251]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[251]_i_2 
       (.I0(\f_permutation_l_/round_in [1028]),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1412]),
        .I4(\out[1585]_i_7_n_0 ),
        .O(\out[251]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[252]_i_1 
       (.I0(\out[252]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[661] ),
        .I2(\out[1443]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[595] ),
        .I4(\out[1238]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [252]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[252]_i_2 
       (.I0(\f_permutation_l_/round_in [1029]),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1413]),
        .I4(\out[1586]_i_7_n_0 ),
        .O(\out[252]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[253]_i_1 
       (.I0(\out[253]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[662] ),
        .I2(\out[1444]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[596] ),
        .I4(\out[1239]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [253]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[253]_i_2 
       (.I0(\f_permutation_l_/round_in [1030]),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1414]),
        .I4(\out[1587]_i_7_n_0 ),
        .O(\out[253]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[254]_i_1 
       (.I0(\out[254]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[663] ),
        .I2(\out[1445]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[597] ),
        .I4(\out[1240]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [254]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[254]_i_2 
       (.I0(\f_permutation_l_/round_in [1031]),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1415]),
        .I4(\out[1588]_i_7_n_0 ),
        .O(\out[254]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[255]_i_1 
       (.I0(\out[255]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[664] ),
        .I2(\out[1446]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[598] ),
        .I4(\out[1241]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [255]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[255]_i_2 
       (.I0(\f_permutation_l_/round_in [1032]),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1416]),
        .I4(\out[1589]_i_7_n_0 ),
        .O(\out[255]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[256]_i_1 
       (.I0(\f_permutation_l_/round_in [1033]),
        .I1(\out[1502]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[665] ),
        .I3(\out[1447]_i_3_n_0 ),
        .I4(\out[256]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [256]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[256]_i_2 
       (.I0(padder_out_1[49]),
        .I1(\f_permutation_l_/out_reg_n_0_[1033] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1033]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[256]_i_3 
       (.I0(\f_permutation_l_/round_in [1410]),
        .I1(\f_permutation_l_/round_in [1345]),
        .I2(\out[1581]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[256]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[257]_i_1 
       (.I0(\f_permutation_l_/round_in [1034]),
        .I1(\out[1503]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[666] ),
        .I3(\out[1448]_i_3_n_0 ),
        .I4(\out[257]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [257]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[257]_i_2 
       (.I0(padder_out_1[50]),
        .I1(\f_permutation_l_/out_reg_n_0_[1034] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1034]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[257]_i_3 
       (.I0(\f_permutation_l_/round_in [1411]),
        .I1(\f_permutation_l_/round_in [1346]),
        .I2(\out[1582]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[257]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[258]_i_1 
       (.I0(\f_permutation_l_/round_in [1035]),
        .I1(\out[1504]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[667] ),
        .I3(\out[1449]_i_3_n_0 ),
        .I4(\out[258]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [258]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[258]_i_2 
       (.I0(padder_out_1[51]),
        .I1(\f_permutation_l_/out_reg_n_0_[1035] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1035]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[258]_i_3 
       (.I0(\f_permutation_l_/round_in [1412]),
        .I1(\f_permutation_l_/round_in [1347]),
        .I2(\out[1583]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[258]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[259]_i_1 
       (.I0(\f_permutation_l_/round_in [1036]),
        .I1(\out[1505]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[668] ),
        .I3(\out[1450]_i_3_n_0 ),
        .I4(\out[259]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [259]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[259]_i_2 
       (.I0(padder_out_1[52]),
        .I1(\f_permutation_l_/out_reg_n_0_[1036] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1036]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[259]_i_3 
       (.I0(\f_permutation_l_/round_in [1413]),
        .I1(\f_permutation_l_/round_in [1348]),
        .I2(\out[1584]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[259]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[25]_i_1 
       (.I0(\out[1539]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[215] ),
        .I2(\out[281]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1058]),
        .I4(\out[1527]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[260]_i_1 
       (.I0(\f_permutation_l_/round_in [1037]),
        .I1(\out[1506]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[669] ),
        .I3(\out[1451]_i_3_n_0 ),
        .I4(\out[260]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [260]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[260]_i_2 
       (.I0(padder_out_1[53]),
        .I1(\f_permutation_l_/out_reg_n_0_[1037] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1037]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[260]_i_3 
       (.I0(\f_permutation_l_/round_in [1414]),
        .I1(\f_permutation_l_/round_in [1349]),
        .I2(\out[1585]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[260]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[261]_i_1 
       (.I0(\f_permutation_l_/round_in [1038]),
        .I1(\out[1507]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[670] ),
        .I3(\out[1452]_i_3_n_0 ),
        .I4(\out[261]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [261]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[261]_i_2 
       (.I0(padder_out_1[54]),
        .I1(\f_permutation_l_/out_reg_n_0_[1038] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1038]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[261]_i_3 
       (.I0(\f_permutation_l_/round_in [1415]),
        .I1(\f_permutation_l_/round_in [1350]),
        .I2(\out[1586]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[261]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[262]_i_1 
       (.I0(\f_permutation_l_/round_in [1039]),
        .I1(\out[1508]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[671] ),
        .I3(\out[1453]_i_3_n_0 ),
        .I4(\out[262]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [262]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[262]_i_2 
       (.I0(padder_out_1[55]),
        .I1(\f_permutation_l_/out_reg_n_0_[1039] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1039]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[262]_i_3 
       (.I0(\f_permutation_l_/round_in [1416]),
        .I1(\f_permutation_l_/round_in [1351]),
        .I2(\out[1587]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[262]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[263]_i_1 
       (.I0(\f_permutation_l_/round_in [1040]),
        .I1(\out[1509]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[672] ),
        .I3(\out[1454]_i_3_n_0 ),
        .I4(\out[263]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [263]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[263]_i_2 
       (.I0(padder_out_1[40]),
        .I1(\f_permutation_l_/out_reg_n_0_[1040] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1040]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[263]_i_3 
       (.I0(\f_permutation_l_/round_in [1417]),
        .I1(\f_permutation_l_/round_in [1352]),
        .I2(\out[1588]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[263]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[264]_i_1 
       (.I0(\f_permutation_l_/round_in [1041]),
        .I1(\out[1510]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[673] ),
        .I3(\out[1455]_i_3_n_0 ),
        .I4(\out[264]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [264]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[264]_i_2 
       (.I0(padder_out_1[41]),
        .I1(\f_permutation_l_/out_reg_n_0_[1041] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1041]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[264]_i_3 
       (.I0(\f_permutation_l_/round_in [1418]),
        .I1(\f_permutation_l_/round_in [1353]),
        .I2(\out[1589]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[264]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[265]_i_1 
       (.I0(\f_permutation_l_/round_in [1042]),
        .I1(\out[1511]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[674] ),
        .I3(\out[1456]_i_3_n_0 ),
        .I4(\out[265]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [265]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[265]_i_2 
       (.I0(padder_out_1[42]),
        .I1(\f_permutation_l_/out_reg_n_0_[1042] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1042]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[265]_i_3 
       (.I0(\f_permutation_l_/round_in [1419]),
        .I1(\f_permutation_l_/round_in [1354]),
        .I2(\out[1590]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[265]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[266]_i_1 
       (.I0(\f_permutation_l_/round_in [1043]),
        .I1(\out[1512]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[675] ),
        .I3(\out[1457]_i_3_n_0 ),
        .I4(\out[266]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [266]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[266]_i_2 
       (.I0(padder_out_1[43]),
        .I1(\f_permutation_l_/out_reg_n_0_[1043] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1043]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[266]_i_3 
       (.I0(\f_permutation_l_/round_in [1420]),
        .I1(\f_permutation_l_/round_in [1355]),
        .I2(\out[1591]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[266]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[267]_i_1 
       (.I0(\f_permutation_l_/round_in [1044]),
        .I1(\out[1513]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[676] ),
        .I3(\out[1458]_i_3_n_0 ),
        .I4(\out[267]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [267]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[267]_i_2 
       (.I0(padder_out_1[44]),
        .I1(\f_permutation_l_/out_reg_n_0_[1044] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1044]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[267]_i_3 
       (.I0(\f_permutation_l_/round_in [1421]),
        .I1(\f_permutation_l_/round_in [1356]),
        .I2(\out[1592]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[267]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[268]_i_1 
       (.I0(\f_permutation_l_/round_in [1045]),
        .I1(\out[1514]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[677] ),
        .I3(\out[1459]_i_3_n_0 ),
        .I4(\out[268]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [268]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[268]_i_2 
       (.I0(padder_out_1[45]),
        .I1(\f_permutation_l_/out_reg_n_0_[1045] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1045]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[268]_i_3 
       (.I0(\f_permutation_l_/round_in [1422]),
        .I1(\f_permutation_l_/round_in [1357]),
        .I2(\out[1593]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[268]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[269]_i_1 
       (.I0(\f_permutation_l_/round_in [1046]),
        .I1(\out[1515]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[678] ),
        .I3(\out[1460]_i_3_n_0 ),
        .I4(\out[269]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [269]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[269]_i_2 
       (.I0(padder_out_1[46]),
        .I1(\f_permutation_l_/out_reg_n_0_[1046] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1046]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[269]_i_3 
       (.I0(\f_permutation_l_/round_in [1423]),
        .I1(\f_permutation_l_/round_in [1358]),
        .I2(\out[1594]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[269]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[26]_i_1 
       (.I0(\out[1540]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[216] ),
        .I2(\out[282]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1059]),
        .I4(\out[1528]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[270]_i_1 
       (.I0(\f_permutation_l_/round_in [1047]),
        .I1(\out[1516]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[679] ),
        .I3(\out[1461]_i_3_n_0 ),
        .I4(\out[270]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [270]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[270]_i_2 
       (.I0(padder_out_1[47]),
        .I1(\f_permutation_l_/out_reg_n_0_[1047] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1047]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[270]_i_3 
       (.I0(\f_permutation_l_/round_in [1424]),
        .I1(\f_permutation_l_/round_in [1359]),
        .I2(\out[1595]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[270]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[271]_i_1 
       (.I0(\f_permutation_l_/round_in [1048]),
        .I1(\out[1517]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[680] ),
        .I3(\out[1462]_i_3_n_0 ),
        .I4(\out[271]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [271]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[271]_i_2 
       (.I0(padder_out_1[32]),
        .I1(\f_permutation_l_/out_reg_n_0_[1048] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1048]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[271]_i_3 
       (.I0(\f_permutation_l_/round_in [1425]),
        .I1(\f_permutation_l_/round_in [1360]),
        .I2(\out[1596]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[271]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[272]_i_1 
       (.I0(\f_permutation_l_/round_in [1049]),
        .I1(\out[1518]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[681] ),
        .I3(\out[1463]_i_3_n_0 ),
        .I4(\out[272]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [272]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[272]_i_2 
       (.I0(padder_out_1[33]),
        .I1(\f_permutation_l_/out_reg_n_0_[1049] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1049]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[272]_i_3 
       (.I0(\f_permutation_l_/round_in [1426]),
        .I1(\f_permutation_l_/round_in [1361]),
        .I2(\out[1597]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[272]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[273]_i_1 
       (.I0(\f_permutation_l_/round_in [1050]),
        .I1(\out[1519]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[682] ),
        .I3(\out[1464]_i_3_n_0 ),
        .I4(\out[273]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [273]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[273]_i_2 
       (.I0(padder_out_1[34]),
        .I1(\f_permutation_l_/out_reg_n_0_[1050] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1050]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[273]_i_3 
       (.I0(\f_permutation_l_/round_in [1427]),
        .I1(\f_permutation_l_/round_in [1362]),
        .I2(\out[1598]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[273]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[274]_i_1 
       (.I0(\f_permutation_l_/round_in [1051]),
        .I1(\out[1520]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[683] ),
        .I3(\out[1465]_i_3_n_0 ),
        .I4(\out[274]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [274]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[274]_i_2 
       (.I0(padder_out_1[35]),
        .I1(\f_permutation_l_/out_reg_n_0_[1051] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1051]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[274]_i_3 
       (.I0(\f_permutation_l_/round_in [1428]),
        .I1(\f_permutation_l_/round_in [1363]),
        .I2(\out[1599]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[274]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[275]_i_1 
       (.I0(\f_permutation_l_/round_in [1052]),
        .I1(\out[1521]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[684] ),
        .I3(\out[1466]_i_3_n_0 ),
        .I4(\out[275]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [275]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[275]_i_2 
       (.I0(padder_out_1[36]),
        .I1(\f_permutation_l_/out_reg_n_0_[1052] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1052]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[275]_i_3 
       (.I0(\f_permutation_l_/round_in [1429]),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1493]),
        .I4(\out[1536]_i_14_n_0 ),
        .O(\out[275]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[276]_i_1 
       (.I0(\f_permutation_l_/round_in [1053]),
        .I1(\out[1522]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[685] ),
        .I3(\out[1467]_i_3_n_0 ),
        .I4(\out[276]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [276]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[276]_i_2 
       (.I0(padder_out_1[37]),
        .I1(\f_permutation_l_/out_reg_n_0_[1053] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1053]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[276]_i_3 
       (.I0(\f_permutation_l_/round_in [1430]),
        .I1(\f_permutation_l_/round_in [1365]),
        .I2(\out[1537]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1494]),
        .I4(\out[1537]_i_10_n_0 ),
        .O(\out[276]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[277]_i_1 
       (.I0(\f_permutation_l_/round_in [1054]),
        .I1(\out[1523]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[686] ),
        .I3(\out[1468]_i_3_n_0 ),
        .I4(\out[277]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [277]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[277]_i_2 
       (.I0(padder_out_1[38]),
        .I1(\f_permutation_l_/out_reg_n_0_[1054] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1054]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[277]_i_3 
       (.I0(\f_permutation_l_/round_in [1431]),
        .I1(\f_permutation_l_/round_in [1366]),
        .I2(\out[1538]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1495]),
        .I4(\out[1538]_i_9_n_0 ),
        .O(\out[277]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[278]_i_1 
       (.I0(\f_permutation_l_/round_in [1055]),
        .I1(\out[1524]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[687] ),
        .I3(\out[1469]_i_3_n_0 ),
        .I4(\out[278]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [278]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[278]_i_2 
       (.I0(padder_out_1[39]),
        .I1(\f_permutation_l_/out_reg_n_0_[1055] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1055]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[278]_i_3 
       (.I0(\f_permutation_l_/round_in [1432]),
        .I1(\out[1539]_i_12_n_0 ),
        .I2(\f_permutation_l_/round_in [1367]),
        .I3(\f_permutation_l_/round_in [1496]),
        .I4(\out[1539]_i_14_n_0 ),
        .O(\out[278]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[279]_i_1 
       (.I0(\f_permutation_l_/round_in [1056]),
        .I1(\out[1525]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[688] ),
        .I3(\out[1470]_i_3_n_0 ),
        .I4(\out[279]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [279]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[279]_i_2 
       (.I0(padder_out_1[24]),
        .I1(\f_permutation_l_/out_reg_n_0_[1056] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1056]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[279]_i_3 
       (.I0(\f_permutation_l_/round_in [1433]),
        .I1(\f_permutation_l_/round_in [1368]),
        .I2(\out[1540]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1497]),
        .I4(\out[1540]_i_9_n_0 ),
        .O(\out[279]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[27]_i_1 
       (.I0(\out[1541]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[217] ),
        .I2(\out[283]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1060]),
        .I4(\out[1529]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[280]_i_1 
       (.I0(\f_permutation_l_/round_in [1057]),
        .I1(\out[1526]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[689] ),
        .I3(\out[1471]_i_3_n_0 ),
        .I4(\out[280]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [280]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[280]_i_2 
       (.I0(padder_out_1[25]),
        .I1(\f_permutation_l_/out_reg_n_0_[1057] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1057]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[280]_i_3 
       (.I0(\f_permutation_l_/round_in [1434]),
        .I1(\f_permutation_l_/round_in [1369]),
        .I2(\out[1541]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1498]),
        .I4(\out[1541]_i_9_n_0 ),
        .O(\out[280]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[281]_i_1 
       (.I0(\f_permutation_l_/round_in [1058]),
        .I1(\out[1527]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[690] ),
        .I3(\out[1408]_i_3_n_0 ),
        .I4(\out[281]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [281]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[281]_i_2 
       (.I0(padder_out_1[26]),
        .I1(\f_permutation_l_/out_reg_n_0_[1058] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1058]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[281]_i_3 
       (.I0(\f_permutation_l_/round_in [1435]),
        .I1(\f_permutation_l_/round_in [1370]),
        .I2(\out[1542]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1499]),
        .I4(\out[1542]_i_11_n_0 ),
        .O(\out[281]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[282]_i_1 
       (.I0(\f_permutation_l_/round_in [1059]),
        .I1(\out[1528]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[691] ),
        .I3(\out[1409]_i_3_n_0 ),
        .I4(\out[282]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [282]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[282]_i_2 
       (.I0(padder_out_1[27]),
        .I1(\f_permutation_l_/out_reg_n_0_[1059] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1059]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[282]_i_3 
       (.I0(\f_permutation_l_/round_in [1436]),
        .I1(\f_permutation_l_/round_in [1371]),
        .I2(\out[1543]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1500]),
        .I4(\out[1543]_i_11_n_0 ),
        .O(\out[282]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[283]_i_1 
       (.I0(\f_permutation_l_/round_in [1060]),
        .I1(\out[1529]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[692] ),
        .I3(\out[1410]_i_3_n_0 ),
        .I4(\out[283]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [283]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[283]_i_2 
       (.I0(padder_out_1[28]),
        .I1(\f_permutation_l_/out_reg_n_0_[1060] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1060]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[283]_i_3 
       (.I0(\f_permutation_l_/round_in [1437]),
        .I1(\f_permutation_l_/round_in [1372]),
        .I2(\out[1544]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1501]),
        .I4(\out[1544]_i_9_n_0 ),
        .O(\out[283]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[284]_i_1 
       (.I0(\f_permutation_l_/round_in [1061]),
        .I1(\out[1530]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[693] ),
        .I3(\out[1411]_i_2_n_0 ),
        .I4(\out[284]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [284]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[284]_i_2 
       (.I0(padder_out_1[29]),
        .I1(\f_permutation_l_/out_reg_n_0_[1061] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1061]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[284]_i_3 
       (.I0(\f_permutation_l_/round_in [1438]),
        .I1(\f_permutation_l_/round_in [1373]),
        .I2(\out[1545]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1502]),
        .I4(\out[1545]_i_9_n_0 ),
        .O(\out[284]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[285]_i_1 
       (.I0(\f_permutation_l_/round_in [1062]),
        .I1(\out[1531]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[694] ),
        .I3(\out[1412]_i_3_n_0 ),
        .I4(\out[285]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [285]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[285]_i_2 
       (.I0(padder_out_1[30]),
        .I1(\f_permutation_l_/out_reg_n_0_[1062] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1062]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[285]_i_3 
       (.I0(\f_permutation_l_/round_in [1439]),
        .I1(\f_permutation_l_/round_in [1374]),
        .I2(\out[1546]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1503]),
        .I4(\out[1546]_i_9_n_0 ),
        .O(\out[285]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[286]_i_1 
       (.I0(\f_permutation_l_/round_in [1063]),
        .I1(\out[1532]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[695] ),
        .I3(\out[1413]_i_3_n_0 ),
        .I4(\out[286]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [286]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[286]_i_2 
       (.I0(padder_out_1[31]),
        .I1(\f_permutation_l_/out_reg_n_0_[1063] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1063]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[286]_i_3 
       (.I0(\f_permutation_l_/round_in [1440]),
        .I1(\f_permutation_l_/round_in [1375]),
        .I2(\out[1547]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1504]),
        .I4(\out[1547]_i_9_n_0 ),
        .O(\out[286]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[287]_i_1 
       (.I0(\f_permutation_l_/round_in [1064]),
        .I1(\out[1533]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[696] ),
        .I3(\out[1414]_i_3_n_0 ),
        .I4(\out[287]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [287]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[287]_i_2 
       (.I0(padder_out_1[16]),
        .I1(\f_permutation_l_/out_reg_n_0_[1064] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1064]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[287]_i_3 
       (.I0(\f_permutation_l_/round_in [1441]),
        .I1(\f_permutation_l_/round_in [1376]),
        .I2(\out[1548]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1505]),
        .I4(\out[1548]_i_9_n_0 ),
        .O(\out[287]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[288]_i_1 
       (.I0(\f_permutation_l_/round_in [1065]),
        .I1(\out[1534]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[697] ),
        .I3(\out[1415]_i_3_n_0 ),
        .I4(\out[288]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [288]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[288]_i_2 
       (.I0(padder_out_1[17]),
        .I1(\f_permutation_l_/out_reg_n_0_[1065] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1065]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[288]_i_3 
       (.I0(\f_permutation_l_/round_in [1442]),
        .I1(\f_permutation_l_/round_in [1377]),
        .I2(\out[1549]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1506]),
        .I4(\out[1549]_i_9_n_0 ),
        .O(\out[288]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[289]_i_1 
       (.I0(\f_permutation_l_/round_in [1066]),
        .I1(\out[1535]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[698] ),
        .I3(\out[1416]_i_3_n_0 ),
        .I4(\out[289]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [289]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[289]_i_2 
       (.I0(padder_out_1[18]),
        .I1(\f_permutation_l_/out_reg_n_0_[1066] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1066]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[289]_i_3 
       (.I0(\f_permutation_l_/round_in [1443]),
        .I1(\f_permutation_l_/round_in [1378]),
        .I2(\out[1550]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1507]),
        .I4(\out[1550]_i_9_n_0 ),
        .O(\out[289]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[28]_i_1 
       (.I0(\out[1542]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[218] ),
        .I2(\out[284]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1061]),
        .I4(\out[1530]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[290]_i_1 
       (.I0(\f_permutation_l_/round_in [1067]),
        .I1(\out[1472]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[699] ),
        .I3(\out[1417]_i_3_n_0 ),
        .I4(\out[290]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [290]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[290]_i_2 
       (.I0(padder_out_1[19]),
        .I1(\f_permutation_l_/out_reg_n_0_[1067] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1067]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[290]_i_3 
       (.I0(\f_permutation_l_/round_in [1444]),
        .I1(\f_permutation_l_/round_in [1379]),
        .I2(\out[1551]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1508]),
        .I4(\out[1551]_i_10_n_0 ),
        .O(\out[290]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[291]_i_1 
       (.I0(\f_permutation_l_/round_in [1068]),
        .I1(\out[1473]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[700] ),
        .I3(\out[1418]_i_3_n_0 ),
        .I4(\out[291]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [291]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[291]_i_2 
       (.I0(padder_out_1[20]),
        .I1(\f_permutation_l_/out_reg_n_0_[1068] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1068]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[291]_i_3 
       (.I0(\f_permutation_l_/round_in [1445]),
        .I1(\f_permutation_l_/round_in [1380]),
        .I2(\out[1552]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1509]),
        .I4(\out[1552]_i_9_n_0 ),
        .O(\out[291]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[292]_i_1 
       (.I0(\f_permutation_l_/round_in [1069]),
        .I1(\out[1474]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[701] ),
        .I3(\out[1419]_i_3_n_0 ),
        .I4(\out[292]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [292]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[292]_i_2 
       (.I0(padder_out_1[21]),
        .I1(\f_permutation_l_/out_reg_n_0_[1069] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1069]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[292]_i_3 
       (.I0(\f_permutation_l_/round_in [1446]),
        .I1(\f_permutation_l_/round_in [1381]),
        .I2(\out[1553]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1510]),
        .I4(\out[1553]_i_9_n_0 ),
        .O(\out[292]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[293]_i_1 
       (.I0(\f_permutation_l_/round_in [1070]),
        .I1(\out[1475]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[702] ),
        .I3(\out[1420]_i_3_n_0 ),
        .I4(\out[293]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [293]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[293]_i_2 
       (.I0(padder_out_1[22]),
        .I1(\f_permutation_l_/out_reg_n_0_[1070] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1070]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[293]_i_3 
       (.I0(\f_permutation_l_/round_in [1447]),
        .I1(\f_permutation_l_/round_in [1382]),
        .I2(\out[1554]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1511]),
        .I4(\out[1554]_i_9_n_0 ),
        .O(\out[293]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[294]_i_1 
       (.I0(\f_permutation_l_/round_in [1071]),
        .I1(\out[1476]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[703] ),
        .I3(\out[1421]_i_3_n_0 ),
        .I4(\out[294]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [294]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[294]_i_2 
       (.I0(padder_out_1[23]),
        .I1(\f_permutation_l_/out_reg_n_0_[1071] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1071]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[294]_i_3 
       (.I0(\f_permutation_l_/round_in [1448]),
        .I1(\f_permutation_l_/round_in [1383]),
        .I2(\out[1555]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1512]),
        .I4(\out[1555]_i_9_n_0 ),
        .O(\out[294]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[295]_i_1 
       (.I0(\f_permutation_l_/round_in [1072]),
        .I1(\out[1477]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[640] ),
        .I3(\out[1422]_i_3_n_0 ),
        .I4(\out[295]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [295]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[295]_i_2 
       (.I0(padder_out_1[8]),
        .I1(\f_permutation_l_/out_reg_n_0_[1072] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1072]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[295]_i_3 
       (.I0(\f_permutation_l_/round_in [1449]),
        .I1(\f_permutation_l_/round_in [1384]),
        .I2(\out[1556]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1513]),
        .I4(\out[1556]_i_10_n_0 ),
        .O(\out[295]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[296]_i_1 
       (.I0(\f_permutation_l_/round_in [1073]),
        .I1(\out[1478]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[641] ),
        .I3(\out[1423]_i_3_n_0 ),
        .I4(\out[296]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [296]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[296]_i_2 
       (.I0(padder_out_1[9]),
        .I1(\f_permutation_l_/out_reg_n_0_[1073] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1073]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[296]_i_3 
       (.I0(\f_permutation_l_/round_in [1450]),
        .I1(\f_permutation_l_/round_in [1385]),
        .I2(\out[1557]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1514]),
        .I4(\out[1557]_i_9_n_0 ),
        .O(\out[296]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[297]_i_1 
       (.I0(\f_permutation_l_/round_in [1074]),
        .I1(\out[1479]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[642] ),
        .I3(\out[1424]_i_3_n_0 ),
        .I4(\out[297]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [297]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[297]_i_2 
       (.I0(padder_out_1[10]),
        .I1(\f_permutation_l_/out_reg_n_0_[1074] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1074]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[297]_i_3 
       (.I0(\f_permutation_l_/round_in [1451]),
        .I1(\f_permutation_l_/round_in [1386]),
        .I2(\out[1558]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1515]),
        .I4(\out[1558]_i_9_n_0 ),
        .O(\out[297]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[298]_i_1 
       (.I0(\f_permutation_l_/round_in [1075]),
        .I1(\out[1480]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[643] ),
        .I3(\out[1425]_i_3_n_0 ),
        .I4(\out[298]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [298]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[298]_i_2 
       (.I0(padder_out_1[11]),
        .I1(\f_permutation_l_/out_reg_n_0_[1075] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1075]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[298]_i_3 
       (.I0(\f_permutation_l_/round_in [1452]),
        .I1(\f_permutation_l_/round_in [1387]),
        .I2(\out[1559]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1516]),
        .I4(\out[1559]_i_9_n_0 ),
        .O(\out[298]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[299]_i_1 
       (.I0(\f_permutation_l_/round_in [1076]),
        .I1(\out[1481]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[644] ),
        .I3(\out[1426]_i_3_n_0 ),
        .I4(\out[299]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [299]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[299]_i_2 
       (.I0(padder_out_1[12]),
        .I1(\f_permutation_l_/out_reg_n_0_[1076] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1076]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[299]_i_3 
       (.I0(\f_permutation_l_/round_in [1453]),
        .I1(\f_permutation_l_/round_in [1388]),
        .I2(\out[1560]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1517]),
        .I4(\out[1560]_i_9_n_0 ),
        .O(\out[299]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[29]_i_1 
       (.I0(\out[1287]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[219] ),
        .I2(\out[285]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1062]),
        .I4(\out[1531]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[2]_i_1 
       (.I0(\out[1580]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[192] ),
        .I2(\out[258]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1035]),
        .I4(\out[1504]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[300]_i_1 
       (.I0(\f_permutation_l_/round_in [1077]),
        .I1(\out[1482]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[645] ),
        .I3(\out[1427]_i_3_n_0 ),
        .I4(\out[300]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [300]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[300]_i_2 
       (.I0(padder_out_1[13]),
        .I1(\f_permutation_l_/out_reg_n_0_[1077] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1077]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[300]_i_3 
       (.I0(\f_permutation_l_/round_in [1454]),
        .I1(\f_permutation_l_/round_in [1389]),
        .I2(\out[1561]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1518]),
        .I4(\out[1561]_i_9_n_0 ),
        .O(\out[300]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[301]_i_1 
       (.I0(\f_permutation_l_/round_in [1078]),
        .I1(\out[1483]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[646] ),
        .I3(\out[1428]_i_3_n_0 ),
        .I4(\out[301]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [301]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[301]_i_2 
       (.I0(padder_out_1[14]),
        .I1(\f_permutation_l_/out_reg_n_0_[1078] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1078]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[301]_i_3 
       (.I0(\f_permutation_l_/round_in [1455]),
        .I1(\f_permutation_l_/round_in [1390]),
        .I2(\out[1562]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1519]),
        .I4(\out[1562]_i_9_n_0 ),
        .O(\out[301]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[302]_i_1 
       (.I0(\f_permutation_l_/round_in [1079]),
        .I1(\out[1484]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[647] ),
        .I3(\out[1429]_i_3_n_0 ),
        .I4(\out[302]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [302]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[302]_i_2 
       (.I0(padder_out_1[15]),
        .I1(\f_permutation_l_/out_reg_n_0_[1079] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1079]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[302]_i_3 
       (.I0(\f_permutation_l_/round_in [1456]),
        .I1(\f_permutation_l_/round_in [1391]),
        .I2(\out[1563]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1520]),
        .I4(\out[1563]_i_9_n_0 ),
        .O(\out[302]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[303]_i_1 
       (.I0(\f_permutation_l_/round_in [1080]),
        .I1(\out[1485]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[648] ),
        .I3(\out[1430]_i_3_n_0 ),
        .I4(\out[303]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [303]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[303]_i_2 
       (.I0(padder_out_1[0]),
        .I1(\f_permutation_l_/out_reg_n_0_[1080] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1080]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[303]_i_3 
       (.I0(\f_permutation_l_/round_in [1457]),
        .I1(\f_permutation_l_/round_in [1392]),
        .I2(\out[1564]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1521]),
        .I4(\out[1564]_i_9_n_0 ),
        .O(\out[303]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[304]_i_1 
       (.I0(\f_permutation_l_/round_in [1081]),
        .I1(\out[1486]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[649] ),
        .I3(\out[1431]_i_3_n_0 ),
        .I4(\out[304]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [304]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[304]_i_2 
       (.I0(padder_out_1[1]),
        .I1(\f_permutation_l_/out_reg_n_0_[1081] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1081]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[304]_i_3 
       (.I0(\f_permutation_l_/round_in [1458]),
        .I1(\f_permutation_l_/round_in [1393]),
        .I2(\out[1565]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1522]),
        .I4(\out[1565]_i_9_n_0 ),
        .O(\out[304]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[305]_i_1 
       (.I0(\f_permutation_l_/round_in [1082]),
        .I1(\out[1487]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[650] ),
        .I3(\out[1432]_i_3_n_0 ),
        .I4(\out[305]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [305]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[305]_i_2 
       (.I0(padder_out_1[2]),
        .I1(\f_permutation_l_/out_reg_n_0_[1082] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1082]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[305]_i_3 
       (.I0(\f_permutation_l_/round_in [1459]),
        .I1(\f_permutation_l_/round_in [1394]),
        .I2(\out[1566]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1523]),
        .I4(\out[1566]_i_9_n_0 ),
        .O(\out[305]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[306]_i_1 
       (.I0(\f_permutation_l_/round_in [1083]),
        .I1(\out[1488]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[651] ),
        .I3(\out[1433]_i_3_n_0 ),
        .I4(\out[306]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [306]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[306]_i_2 
       (.I0(padder_out_1[3]),
        .I1(\f_permutation_l_/out_reg_n_0_[1083] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1083]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[306]_i_3 
       (.I0(\f_permutation_l_/round_in [1460]),
        .I1(\f_permutation_l_/round_in [1395]),
        .I2(\out[1567]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1524]),
        .I4(\out[1567]_i_10_n_0 ),
        .O(\out[306]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[307]_i_1 
       (.I0(\f_permutation_l_/round_in [1084]),
        .I1(\out[1489]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[652] ),
        .I3(\out[1434]_i_3_n_0 ),
        .I4(\out[307]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [307]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[307]_i_2 
       (.I0(padder_out_1[4]),
        .I1(\f_permutation_l_/out_reg_n_0_[1084] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1084]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[307]_i_3 
       (.I0(\f_permutation_l_/round_in [1461]),
        .I1(\f_permutation_l_/round_in [1396]),
        .I2(\out[1568]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1525]),
        .I4(\out[1568]_i_9_n_0 ),
        .O(\out[307]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[308]_i_1 
       (.I0(\f_permutation_l_/round_in [1085]),
        .I1(\out[1490]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[653] ),
        .I3(\out[1435]_i_3_n_0 ),
        .I4(\out[308]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [308]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[308]_i_2 
       (.I0(padder_out_1[5]),
        .I1(\f_permutation_l_/out_reg_n_0_[1085] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1085]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[308]_i_3 
       (.I0(\f_permutation_l_/round_in [1462]),
        .I1(\f_permutation_l_/round_in [1397]),
        .I2(\out[1569]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1526]),
        .I4(\out[1569]_i_9_n_0 ),
        .O(\out[308]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[309]_i_1 
       (.I0(\f_permutation_l_/round_in [1086]),
        .I1(\out[1491]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[654] ),
        .I3(\out[1436]_i_3_n_0 ),
        .I4(\out[309]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [309]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[309]_i_2 
       (.I0(padder_out_1[6]),
        .I1(\f_permutation_l_/out_reg_n_0_[1086] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1086]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[309]_i_3 
       (.I0(\f_permutation_l_/round_in [1463]),
        .I1(\f_permutation_l_/round_in [1398]),
        .I2(\out[1570]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1527]),
        .I4(\out[1570]_i_9_n_0 ),
        .O(\out[309]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[30]_i_1 
       (.I0(\out[1544]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[220] ),
        .I2(\out[286]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1063]),
        .I4(\out[1532]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[310]_i_1 
       (.I0(\f_permutation_l_/round_in [1087]),
        .I1(\out[1492]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[655] ),
        .I3(\out[1437]_i_3_n_0 ),
        .I4(\out[310]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [310]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[310]_i_2 
       (.I0(padder_out_1[7]),
        .I1(\f_permutation_l_/out_reg_n_0_[1087] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1087]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[310]_i_3 
       (.I0(\f_permutation_l_/round_in [1464]),
        .I1(\f_permutation_l_/round_in [1399]),
        .I2(\out[1571]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1528]),
        .I4(\out[1571]_i_9_n_0 ),
        .O(\out[310]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[311]_i_1 
       (.I0(\f_permutation_l_/round_in [1024]),
        .I1(\out[1493]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[656] ),
        .I3(\out[1438]_i_3_n_0 ),
        .I4(\out[311]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [311]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[311]_i_2 
       (.I0(padder_out_1[56]),
        .I1(\f_permutation_l_/out_reg_n_0_[1024] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1024]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[311]_i_3 
       (.I0(\f_permutation_l_/round_in [1465]),
        .I1(\f_permutation_l_/round_in [1400]),
        .I2(\out[1572]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1529]),
        .I4(\out[1572]_i_9_n_0 ),
        .O(\out[311]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[312]_i_1 
       (.I0(\f_permutation_l_/round_in [1025]),
        .I1(\out[1494]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[657] ),
        .I3(\out[1439]_i_3_n_0 ),
        .I4(\out[312]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [312]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[312]_i_2 
       (.I0(padder_out_1[57]),
        .I1(\f_permutation_l_/out_reg_n_0_[1025] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1025]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[312]_i_3 
       (.I0(\f_permutation_l_/round_in [1466]),
        .I1(\f_permutation_l_/round_in [1401]),
        .I2(\out[1573]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1530]),
        .I4(\out[1573]_i_9_n_0 ),
        .O(\out[312]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[313]_i_1 
       (.I0(\f_permutation_l_/round_in [1026]),
        .I1(\out[1495]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[658] ),
        .I3(\out[1440]_i_3_n_0 ),
        .I4(\out[313]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [313]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[313]_i_2 
       (.I0(padder_out_1[58]),
        .I1(\f_permutation_l_/out_reg_n_0_[1026] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1026]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[313]_i_3 
       (.I0(\f_permutation_l_/round_in [1467]),
        .I1(\f_permutation_l_/round_in [1402]),
        .I2(\out[1574]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1531]),
        .I4(\out[1574]_i_9_n_0 ),
        .O(\out[313]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[314]_i_1 
       (.I0(\f_permutation_l_/round_in [1027]),
        .I1(\out[1496]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[659] ),
        .I3(\out[1441]_i_3_n_0 ),
        .I4(\out[314]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [314]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[314]_i_2 
       (.I0(padder_out_1[59]),
        .I1(\f_permutation_l_/out_reg_n_0_[1027] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1027]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[314]_i_3 
       (.I0(\f_permutation_l_/round_in [1468]),
        .I1(\f_permutation_l_/round_in [1403]),
        .I2(\out[1575]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1532]),
        .I4(\out[1575]_i_9_n_0 ),
        .O(\out[314]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[315]_i_1 
       (.I0(\f_permutation_l_/round_in [1028]),
        .I1(\out[1497]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[660] ),
        .I3(\out[1442]_i_3_n_0 ),
        .I4(\out[315]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [315]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[315]_i_2 
       (.I0(padder_out_1[60]),
        .I1(\f_permutation_l_/out_reg_n_0_[1028] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1028]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[315]_i_3 
       (.I0(\f_permutation_l_/round_in [1469]),
        .I1(\f_permutation_l_/round_in [1404]),
        .I2(\out[1576]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1533]),
        .I4(\out[1576]_i_9_n_0 ),
        .O(\out[315]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[316]_i_1 
       (.I0(\f_permutation_l_/round_in [1029]),
        .I1(\out[1498]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[661] ),
        .I3(\out[1443]_i_3_n_0 ),
        .I4(\out[316]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [316]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[316]_i_2 
       (.I0(padder_out_1[61]),
        .I1(\f_permutation_l_/out_reg_n_0_[1029] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1029]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[316]_i_3 
       (.I0(\f_permutation_l_/round_in [1470]),
        .I1(\f_permutation_l_/round_in [1405]),
        .I2(\out[1577]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1534]),
        .I4(\out[1577]_i_9_n_0 ),
        .O(\out[316]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[317]_i_1 
       (.I0(\f_permutation_l_/round_in [1030]),
        .I1(\out[1499]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[662] ),
        .I3(\out[1444]_i_3_n_0 ),
        .I4(\out[317]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [317]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[317]_i_2 
       (.I0(padder_out_1[62]),
        .I1(\f_permutation_l_/out_reg_n_0_[1030] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1030]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[317]_i_3 
       (.I0(\f_permutation_l_/round_in [1471]),
        .I1(\f_permutation_l_/round_in [1406]),
        .I2(\out[1578]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[317]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[318]_i_1 
       (.I0(\f_permutation_l_/round_in [1031]),
        .I1(\out[1500]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[663] ),
        .I3(\out[1445]_i_3_n_0 ),
        .I4(\out[318]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [318]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[318]_i_2 
       (.I0(padder_out_1[63]),
        .I1(\f_permutation_l_/out_reg_n_0_[1031] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1031]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[318]_i_3 
       (.I0(\f_permutation_l_/round_in [1408]),
        .I1(\f_permutation_l_/round_in [1407]),
        .I2(\out[1579]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[318]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[319]_i_1 
       (.I0(\f_permutation_l_/round_in [1032]),
        .I1(\out[1501]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[664] ),
        .I3(\out[1446]_i_3_n_0 ),
        .I4(\out[319]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [319]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[319]_i_2 
       (.I0(padder_out_1[48]),
        .I1(\f_permutation_l_/out_reg_n_0_[1032] ),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1032]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[319]_i_3 
       (.I0(\f_permutation_l_/round_in [1409]),
        .I1(\f_permutation_l_/round_in [1344]),
        .I2(\out[1580]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[319]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[31]_i_1 
       (.I0(\out[1545]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[221] ),
        .I2(\out[287]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1064]),
        .I4(\out[1533]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[320]_i_1 
       (.I0(\out[1501]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[72] ),
        .I2(\out[576]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1244]),
        .I4(\out[1247]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [320]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[321]_i_1 
       (.I0(\out[1502]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[73] ),
        .I2(\out[577]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1245]),
        .I4(\out[1248]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [321]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[322]_i_1 
       (.I0(\out[1503]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[74] ),
        .I2(\out[578]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1246]),
        .I4(\out[1249]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [322]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[323]_i_1 
       (.I0(\out[1504]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[75] ),
        .I2(\out[579]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1247]),
        .I4(\out[1250]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [323]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[324]_i_1 
       (.I0(\out[1505]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[76] ),
        .I2(\out[580]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1248]),
        .I4(\out[1251]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [324]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[325]_i_1 
       (.I0(\out[1506]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[77] ),
        .I2(\out[581]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1249]),
        .I4(\out[1252]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [325]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[326]_i_1 
       (.I0(\out[1507]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[78] ),
        .I2(\out[582]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1250]),
        .I4(\out[1253]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [326]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[327]_i_1 
       (.I0(\out[1508]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[79] ),
        .I2(\out[583]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1251]),
        .I4(\out[1254]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [327]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[328]_i_1 
       (.I0(\out[1509]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[80] ),
        .I2(\out[584]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1252]),
        .I4(\out[1255]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [328]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[329]_i_1 
       (.I0(\out[1510]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[81] ),
        .I2(\out[585]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1253]),
        .I4(\out[1256]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [329]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[32]_i_1 
       (.I0(\out[1546]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[222] ),
        .I2(\out[288]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1065]),
        .I4(\out[1534]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[330]_i_1 
       (.I0(\out[1511]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[82] ),
        .I2(\out[586]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1254]),
        .I4(\out[1257]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [330]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[331]_i_1 
       (.I0(\out[1512]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[83] ),
        .I2(\out[587]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1255]),
        .I4(\out[1258]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [331]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[332]_i_1 
       (.I0(\out[1513]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[84] ),
        .I2(\out[588]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1256]),
        .I4(\out[1259]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [332]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[333]_i_1 
       (.I0(\out[1514]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[85] ),
        .I2(\out[589]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1257]),
        .I4(\out[1260]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [333]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[334]_i_1 
       (.I0(\out[1515]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[86] ),
        .I2(\out[590]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1258]),
        .I4(\out[1261]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [334]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[335]_i_1 
       (.I0(\out[1516]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[87] ),
        .I2(\out[591]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1259]),
        .I4(\out[1262]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [335]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[336]_i_1 
       (.I0(\out[1517]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[88] ),
        .I2(\out[592]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1260]),
        .I4(\out[1263]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [336]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[337]_i_1 
       (.I0(\out[1518]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[89] ),
        .I2(\out[593]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1261]),
        .I4(\out[1264]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [337]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[338]_i_1 
       (.I0(\out[1519]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[90] ),
        .I2(\out[594]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1262]),
        .I4(\out[1265]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [338]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[339]_i_1 
       (.I0(\out[1520]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[91] ),
        .I2(\out[595]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1263]),
        .I4(\out[1266]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [339]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[33]_i_1 
       (.I0(\out[1547]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[223] ),
        .I2(\out[289]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1066]),
        .I4(\out[1535]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[340]_i_1 
       (.I0(\out[1521]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[92] ),
        .I2(\out[596]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1264]),
        .I4(\out[1267]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [340]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[341]_i_1 
       (.I0(\out[1522]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[93] ),
        .I2(\out[597]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1265]),
        .I4(\out[1268]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [341]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[342]_i_1 
       (.I0(\out[1523]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[94] ),
        .I2(\out[598]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1266]),
        .I4(\out[1269]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [342]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[343]_i_1 
       (.I0(\out[1524]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[95] ),
        .I2(\out[599]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1267]),
        .I4(\out[1270]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [343]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[344]_i_1 
       (.I0(\out[1525]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[96] ),
        .I2(\out[600]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1268]),
        .I4(\out[1271]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [344]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[345]_i_1 
       (.I0(\out[1526]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[97] ),
        .I2(\out[601]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1269]),
        .I4(\out[1272]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [345]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[346]_i_1 
       (.I0(\out[1527]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[98] ),
        .I2(\out[602]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1270]),
        .I4(\out[1273]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [346]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[347]_i_1 
       (.I0(\out[1528]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[99] ),
        .I2(\out[603]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1271]),
        .I4(\out[1274]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [347]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[348]_i_1 
       (.I0(\out[1529]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[100] ),
        .I2(\out[604]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1272]),
        .I4(\out[1275]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [348]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[349]_i_1 
       (.I0(\out[1530]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[101] ),
        .I2(\out[605]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1273]),
        .I4(\out[1276]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [349]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[34]_i_1 
       (.I0(\out[1548]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[224] ),
        .I2(\out[290]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1067]),
        .I4(\out[1472]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[350]_i_1 
       (.I0(\out[1531]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[102] ),
        .I2(\out[606]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1274]),
        .I4(\out[1277]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [350]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[351]_i_1 
       (.I0(\out[1532]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[103] ),
        .I2(\out[607]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1275]),
        .I4(\out[1278]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [351]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[352]_i_1 
       (.I0(\out[1533]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[104] ),
        .I2(\out[608]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1276]),
        .I4(\out[1279]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [352]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[353]_i_1 
       (.I0(\out[1534]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[105] ),
        .I2(\out[609]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1277]),
        .I4(\out[1216]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [353]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[354]_i_1 
       (.I0(\out[1535]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[106] ),
        .I2(\out[610]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1278]),
        .I4(\out[1217]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [354]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[355]_i_1 
       (.I0(\out[1472]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[107] ),
        .I2(\out[611]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1279]),
        .I4(\out[1218]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [355]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[356]_i_1 
       (.I0(\out[1473]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[108] ),
        .I2(\out[612]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1216]),
        .I4(\out[1219]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [356]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[357]_i_1 
       (.I0(\out[1474]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[109] ),
        .I2(\out[613]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1217]),
        .I4(\out[1220]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [357]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[358]_i_1 
       (.I0(\out[1475]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[110] ),
        .I2(\out[614]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1218]),
        .I4(\out[1221]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [358]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[359]_i_1 
       (.I0(\out[1476]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[111] ),
        .I2(\out[615]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1219]),
        .I4(\out[1539]_i_6_n_0 ),
        .O(\f_permutation_l_/round_out [359]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[35]_i_1 
       (.I0(\out[1549]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[225] ),
        .I2(\out[291]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1068]),
        .I4(\out[1473]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[360]_i_1 
       (.I0(\out[1477]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[112] ),
        .I2(\out[616]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1220]),
        .I4(\out[1223]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [360]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[361]_i_1 
       (.I0(\out[1478]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[113] ),
        .I2(\out[617]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1221]),
        .I4(\out[1224]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [361]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[362]_i_1 
       (.I0(\out[1479]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[114] ),
        .I2(\out[618]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1222]),
        .I4(\out[1225]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [362]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[363]_i_1 
       (.I0(\out[1480]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[115] ),
        .I2(\out[619]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1223]),
        .I4(\out[1226]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [363]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[364]_i_1 
       (.I0(\out[1481]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[116] ),
        .I2(\out[620]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1224]),
        .I4(\out[1227]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [364]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[365]_i_1 
       (.I0(\out[1482]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[117] ),
        .I2(\out[621]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1225]),
        .I4(\out[1228]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [365]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[366]_i_1 
       (.I0(\out[1483]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[118] ),
        .I2(\out[622]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1226]),
        .I4(\out[1229]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [366]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[367]_i_1 
       (.I0(\out[1484]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[119] ),
        .I2(\out[623]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1227]),
        .I4(\out[1230]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [367]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[368]_i_1 
       (.I0(\out[1485]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[120] ),
        .I2(\out[624]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1228]),
        .I4(\out[1231]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [368]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[369]_i_1 
       (.I0(\out[1486]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[121] ),
        .I2(\out[625]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1229]),
        .I4(\out[1232]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [369]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[36]_i_1 
       (.I0(\out[1550]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[226] ),
        .I2(\out[292]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1069]),
        .I4(\out[1474]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[370]_i_1 
       (.I0(\out[1487]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[122] ),
        .I2(\out[626]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1230]),
        .I4(\out[1233]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [370]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[371]_i_1 
       (.I0(\out[1488]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[123] ),
        .I2(\out[627]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1231]),
        .I4(\out[1234]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [371]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[372]_i_1 
       (.I0(\out[1489]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[124] ),
        .I2(\out[628]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1232]),
        .I4(\out[1235]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [372]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[373]_i_1 
       (.I0(\out[1490]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[125] ),
        .I2(\out[629]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1233]),
        .I4(\out[1236]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [373]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[374]_i_1 
       (.I0(\out[1491]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[126] ),
        .I2(\out[630]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1234]),
        .I4(\out[1237]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [374]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[375]_i_1 
       (.I0(\out[1492]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[127] ),
        .I2(\out[631]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1235]),
        .I4(\out[1238]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [375]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[376]_i_1 
       (.I0(\out[1493]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[64] ),
        .I2(\out[632]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1236]),
        .I4(\out[1239]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [376]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[377]_i_1 
       (.I0(\out[1494]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[65] ),
        .I2(\out[633]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1237]),
        .I4(\out[1240]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [377]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[378]_i_1 
       (.I0(\out[1495]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[66] ),
        .I2(\out[634]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1238]),
        .I4(\out[1241]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [378]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[379]_i_1 
       (.I0(\out[1496]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[67] ),
        .I2(\out[635]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1239]),
        .I4(\out[1242]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [379]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[37]_i_1 
       (.I0(\out[1295]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[227] ),
        .I2(\out[293]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1070]),
        .I4(\out[1475]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[380]_i_1 
       (.I0(\out[1497]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[68] ),
        .I2(\out[636]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1240]),
        .I4(\out[1243]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [380]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[381]_i_1 
       (.I0(\out[1498]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[69] ),
        .I2(\out[637]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1241]),
        .I4(\out[1244]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [381]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[382]_i_1 
       (.I0(\out[1499]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[70] ),
        .I2(\out[638]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1242]),
        .I4(\out[1245]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [382]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[383]_i_1 
       (.I0(\out[1500]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[71] ),
        .I2(\out[639]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1243]),
        .I4(\out[1246]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [383]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[384]_i_1 
       (.I0(\out[1564]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[497] ),
        .I2(\f_permutation_l_/out_reg_n_0_[72] ),
        .I3(\out[1501]_i_3_n_0 ),
        .I4(\out[576]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [384]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[385]_i_1 
       (.I0(\out[1565]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[498] ),
        .I2(\f_permutation_l_/out_reg_n_0_[73] ),
        .I3(\out[1502]_i_3_n_0 ),
        .I4(\out[577]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [385]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[386]_i_1 
       (.I0(\out[1566]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[499] ),
        .I2(\f_permutation_l_/out_reg_n_0_[74] ),
        .I3(\out[1503]_i_2_n_0 ),
        .I4(\out[578]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [386]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[387]_i_1 
       (.I0(\out[1567]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[500] ),
        .I2(\f_permutation_l_/out_reg_n_0_[75] ),
        .I3(\out[1504]_i_3_n_0 ),
        .I4(\out[579]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [387]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[388]_i_1 
       (.I0(\out[1568]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[501] ),
        .I2(\f_permutation_l_/out_reg_n_0_[76] ),
        .I3(\out[1505]_i_3_n_0 ),
        .I4(\out[580]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [388]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[389]_i_1 
       (.I0(\out[1569]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[502] ),
        .I2(\f_permutation_l_/out_reg_n_0_[77] ),
        .I3(\out[1506]_i_3_n_0 ),
        .I4(\out[581]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [389]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[38]_i_1 
       (.I0(\out[1552]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[228] ),
        .I2(\out[294]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1071]),
        .I4(\out[1476]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[390]_i_1 
       (.I0(\out[1570]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[503] ),
        .I2(\f_permutation_l_/out_reg_n_0_[78] ),
        .I3(\out[1507]_i_3_n_0 ),
        .I4(\out[582]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [390]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[391]_i_1 
       (.I0(\out[1571]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[504] ),
        .I2(\f_permutation_l_/out_reg_n_0_[79] ),
        .I3(\out[1508]_i_3_n_0 ),
        .I4(\out[583]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [391]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[392]_i_1 
       (.I0(\out[1572]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[505] ),
        .I2(\f_permutation_l_/out_reg_n_0_[80] ),
        .I3(\out[1509]_i_3_n_0 ),
        .I4(\out[584]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [392]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[393]_i_1 
       (.I0(\out[1573]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[506] ),
        .I2(\f_permutation_l_/out_reg_n_0_[81] ),
        .I3(\out[1510]_i_3_n_0 ),
        .I4(\out[585]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [393]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[394]_i_1 
       (.I0(\out[1574]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[507] ),
        .I2(\f_permutation_l_/out_reg_n_0_[82] ),
        .I3(\out[1511]_i_3_n_0 ),
        .I4(\out[586]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [394]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[395]_i_1 
       (.I0(\out[1575]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[508] ),
        .I2(\f_permutation_l_/out_reg_n_0_[83] ),
        .I3(\out[1512]_i_3_n_0 ),
        .I4(\out[587]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [395]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[396]_i_1 
       (.I0(\out[1576]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[509] ),
        .I2(\f_permutation_l_/out_reg_n_0_[84] ),
        .I3(\out[1513]_i_3_n_0 ),
        .I4(\out[588]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [396]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[397]_i_1 
       (.I0(\out[1577]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[510] ),
        .I2(\f_permutation_l_/out_reg_n_0_[85] ),
        .I3(\out[1514]_i_3_n_0 ),
        .I4(\out[589]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [397]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[398]_i_1 
       (.I0(\out[1578]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[511] ),
        .I2(\f_permutation_l_/out_reg_n_0_[86] ),
        .I3(\out[1515]_i_3_n_0 ),
        .I4(\out[590]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [398]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[399]_i_1 
       (.I0(\out[1579]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[448] ),
        .I2(\f_permutation_l_/out_reg_n_0_[87] ),
        .I3(\out[1516]_i_3_n_0 ),
        .I4(\out[591]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [399]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[39]_i_1 
       (.I0(\out[1553]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[229] ),
        .I2(\out[295]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1072]),
        .I4(\out[1477]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[3]_i_1 
       (.I0(\out[1581]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[193] ),
        .I2(\out[259]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1036]),
        .I4(\out[1505]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[400]_i_1 
       (.I0(\out[1580]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[449] ),
        .I2(\f_permutation_l_/out_reg_n_0_[88] ),
        .I3(\out[1517]_i_3_n_0 ),
        .I4(\out[592]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [400]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[401]_i_1 
       (.I0(\out[1581]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[450] ),
        .I2(\f_permutation_l_/out_reg_n_0_[89] ),
        .I3(\out[1518]_i_3_n_0 ),
        .I4(\out[593]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [401]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[402]_i_1 
       (.I0(\out[1582]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[451] ),
        .I2(\f_permutation_l_/out_reg_n_0_[90] ),
        .I3(\out[1519]_i_3_n_0 ),
        .I4(\out[594]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [402]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[403]_i_1 
       (.I0(\out[1583]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[452] ),
        .I2(\f_permutation_l_/out_reg_n_0_[91] ),
        .I3(\out[1520]_i_3_n_0 ),
        .I4(\out[595]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [403]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[404]_i_1 
       (.I0(\out[1584]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[453] ),
        .I2(\f_permutation_l_/out_reg_n_0_[92] ),
        .I3(\out[1521]_i_3_n_0 ),
        .I4(\out[596]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [404]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[405]_i_1 
       (.I0(\out[1585]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[454] ),
        .I2(\f_permutation_l_/out_reg_n_0_[93] ),
        .I3(\out[1522]_i_3_n_0 ),
        .I4(\out[597]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [405]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[406]_i_1 
       (.I0(\out[1586]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[455] ),
        .I2(\f_permutation_l_/out_reg_n_0_[94] ),
        .I3(\out[1523]_i_3_n_0 ),
        .I4(\out[598]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [406]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[407]_i_1 
       (.I0(\out[1587]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[456] ),
        .I2(\f_permutation_l_/out_reg_n_0_[95] ),
        .I3(\out[1524]_i_3_n_0 ),
        .I4(\out[599]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [407]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[408]_i_1 
       (.I0(\out[1588]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[457] ),
        .I2(\f_permutation_l_/out_reg_n_0_[96] ),
        .I3(\out[1525]_i_3_n_0 ),
        .I4(\out[600]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [408]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[409]_i_1 
       (.I0(\out[1589]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[458] ),
        .I2(\f_permutation_l_/out_reg_n_0_[97] ),
        .I3(\out[1526]_i_3_n_0 ),
        .I4(\out[601]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [409]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[40]_i_1 
       (.I0(\out[1554]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[230] ),
        .I2(\out[296]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1073]),
        .I4(\out[1478]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[410]_i_1 
       (.I0(\out[1590]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[459] ),
        .I2(\f_permutation_l_/out_reg_n_0_[98] ),
        .I3(\out[1527]_i_3_n_0 ),
        .I4(\out[602]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [410]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[411]_i_1 
       (.I0(\out[1591]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[460] ),
        .I2(\f_permutation_l_/out_reg_n_0_[99] ),
        .I3(\out[1528]_i_3_n_0 ),
        .I4(\out[603]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [411]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[412]_i_1 
       (.I0(\out[1592]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[461] ),
        .I2(\f_permutation_l_/out_reg_n_0_[100] ),
        .I3(\out[1529]_i_3_n_0 ),
        .I4(\out[604]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [412]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[413]_i_1 
       (.I0(\out[1593]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[462] ),
        .I2(\f_permutation_l_/out_reg_n_0_[101] ),
        .I3(\out[1530]_i_3_n_0 ),
        .I4(\out[605]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [413]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[414]_i_1 
       (.I0(\out[1594]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[463] ),
        .I2(\f_permutation_l_/out_reg_n_0_[102] ),
        .I3(\out[1531]_i_3_n_0 ),
        .I4(\out[606]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [414]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[415]_i_1 
       (.I0(\out[1595]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[464] ),
        .I2(\f_permutation_l_/out_reg_n_0_[103] ),
        .I3(\out[1532]_i_3_n_0 ),
        .I4(\out[607]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [415]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[416]_i_1 
       (.I0(\out[1596]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[465] ),
        .I2(\f_permutation_l_/out_reg_n_0_[104] ),
        .I3(\out[1533]_i_3_n_0 ),
        .I4(\out[608]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [416]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[417]_i_1 
       (.I0(\out[1597]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[466] ),
        .I2(\f_permutation_l_/out_reg_n_0_[105] ),
        .I3(\out[1534]_i_3_n_0 ),
        .I4(\out[609]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [417]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[418]_i_1 
       (.I0(\out[1598]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[467] ),
        .I2(\f_permutation_l_/out_reg_n_0_[106] ),
        .I3(\out[1535]_i_2_n_0 ),
        .I4(\out[610]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [418]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[419]_i_1 
       (.I0(\out[1599]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[468] ),
        .I2(\f_permutation_l_/out_reg_n_0_[107] ),
        .I3(\out[1472]_i_3_n_0 ),
        .I4(\out[611]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [419]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[41]_i_1 
       (.I0(\out[1555]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[231] ),
        .I2(\out[297]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1074]),
        .I4(\out[1479]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[420]_i_1 
       (.I0(\out[1472]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[469] ),
        .I2(\f_permutation_l_/out_reg_n_0_[108] ),
        .I3(\out[1473]_i_2_n_0 ),
        .I4(\out[612]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [420]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[421]_i_1 
       (.I0(\out[1537]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[470] ),
        .I2(\f_permutation_l_/out_reg_n_0_[109] ),
        .I3(\out[1474]_i_3_n_0 ),
        .I4(\out[613]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [421]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[422]_i_1 
       (.I0(\out[1538]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[471] ),
        .I2(\f_permutation_l_/out_reg_n_0_[110] ),
        .I3(\out[1475]_i_2_n_0 ),
        .I4(\out[614]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [422]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[423]_i_1 
       (.I0(\out[1045]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[472] ),
        .I2(\f_permutation_l_/out_reg_n_0_[111] ),
        .I3(\out[1476]_i_3_n_0 ),
        .I4(\out[615]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [423]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[424]_i_1 
       (.I0(\out[1540]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[473] ),
        .I2(\f_permutation_l_/out_reg_n_0_[112] ),
        .I3(\out[1477]_i_3_n_0 ),
        .I4(\out[616]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [424]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[425]_i_1 
       (.I0(\out[1541]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[474] ),
        .I2(\f_permutation_l_/out_reg_n_0_[113] ),
        .I3(\out[1478]_i_3_n_0 ),
        .I4(\out[617]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [425]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[426]_i_1 
       (.I0(\out[1542]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[475] ),
        .I2(\f_permutation_l_/out_reg_n_0_[114] ),
        .I3(\out[1479]_i_2_n_0 ),
        .I4(\out[618]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [426]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[427]_i_1 
       (.I0(\out[1543]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[476] ),
        .I2(\f_permutation_l_/out_reg_n_0_[115] ),
        .I3(\out[1480]_i_3_n_0 ),
        .I4(\out[619]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [427]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[428]_i_1 
       (.I0(\out[1544]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[477] ),
        .I2(\f_permutation_l_/out_reg_n_0_[116] ),
        .I3(\out[1481]_i_3_n_0 ),
        .I4(\out[620]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [428]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[429]_i_1 
       (.I0(\out[1545]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[478] ),
        .I2(\f_permutation_l_/out_reg_n_0_[117] ),
        .I3(\out[1482]_i_3_n_0 ),
        .I4(\out[621]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [429]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[42]_i_1 
       (.I0(\out[1556]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[232] ),
        .I2(\out[298]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1075]),
        .I4(\out[1480]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[430]_i_1 
       (.I0(\out[1546]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[479] ),
        .I2(\f_permutation_l_/out_reg_n_0_[118] ),
        .I3(\out[1483]_i_3_n_0 ),
        .I4(\out[622]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [430]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[431]_i_1 
       (.I0(\out[1547]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[480] ),
        .I2(\f_permutation_l_/out_reg_n_0_[119] ),
        .I3(\out[1484]_i_3_n_0 ),
        .I4(\out[623]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [431]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[432]_i_1 
       (.I0(\out[1548]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[481] ),
        .I2(\f_permutation_l_/out_reg_n_0_[120] ),
        .I3(\out[1485]_i_3_n_0 ),
        .I4(\out[624]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [432]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[433]_i_1 
       (.I0(\out[1549]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[482] ),
        .I2(\f_permutation_l_/out_reg_n_0_[121] ),
        .I3(\out[1486]_i_3_n_0 ),
        .I4(\out[625]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [433]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[434]_i_1 
       (.I0(\out[1550]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[483] ),
        .I2(\f_permutation_l_/out_reg_n_0_[122] ),
        .I3(\out[1487]_i_2_n_0 ),
        .I4(\out[626]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [434]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[435]_i_1 
       (.I0(\out[1551]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[484] ),
        .I2(\f_permutation_l_/out_reg_n_0_[123] ),
        .I3(\out[1488]_i_3_n_0 ),
        .I4(\out[627]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [435]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[436]_i_1 
       (.I0(\out[1552]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[485] ),
        .I2(\f_permutation_l_/out_reg_n_0_[124] ),
        .I3(\out[1489]_i_3_n_0 ),
        .I4(\out[628]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [436]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[437]_i_1 
       (.I0(\out[1553]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[486] ),
        .I2(\f_permutation_l_/out_reg_n_0_[125] ),
        .I3(\out[1490]_i_3_n_0 ),
        .I4(\out[629]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [437]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[438]_i_1 
       (.I0(\out[1554]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[487] ),
        .I2(\f_permutation_l_/out_reg_n_0_[126] ),
        .I3(\out[1491]_i_3_n_0 ),
        .I4(\out[630]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [438]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[439]_i_1 
       (.I0(\out[1555]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[488] ),
        .I2(\f_permutation_l_/out_reg_n_0_[127] ),
        .I3(\out[1492]_i_3_n_0 ),
        .I4(\out[631]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [439]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[43]_i_1 
       (.I0(\out[1557]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[233] ),
        .I2(\out[299]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1076]),
        .I4(\out[1481]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[440]_i_1 
       (.I0(\out[1556]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[489] ),
        .I2(\f_permutation_l_/out_reg_n_0_[64] ),
        .I3(\out[1493]_i_3_n_0 ),
        .I4(\out[632]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [440]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[441]_i_1 
       (.I0(\out[1557]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[490] ),
        .I2(\f_permutation_l_/out_reg_n_0_[65] ),
        .I3(\out[1494]_i_3_n_0 ),
        .I4(\out[633]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [441]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[442]_i_1 
       (.I0(\out[1558]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[491] ),
        .I2(\f_permutation_l_/out_reg_n_0_[66] ),
        .I3(\out[1495]_i_3_n_0 ),
        .I4(\out[634]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [442]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[443]_i_1 
       (.I0(\out[1559]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[492] ),
        .I2(\f_permutation_l_/out_reg_n_0_[67] ),
        .I3(\out[1496]_i_3_n_0 ),
        .I4(\out[635]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [443]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[444]_i_1 
       (.I0(\out[1560]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[493] ),
        .I2(\f_permutation_l_/out_reg_n_0_[68] ),
        .I3(\out[1497]_i_3_n_0 ),
        .I4(\out[636]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [444]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[445]_i_1 
       (.I0(\out[1561]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[494] ),
        .I2(\f_permutation_l_/out_reg_n_0_[69] ),
        .I3(\out[1498]_i_3_n_0 ),
        .I4(\out[637]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [445]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[446]_i_1 
       (.I0(\out[1562]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[495] ),
        .I2(\f_permutation_l_/out_reg_n_0_[70] ),
        .I3(\out[1499]_i_3_n_0 ),
        .I4(\out[638]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [446]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[447]_i_1 
       (.I0(\out[1563]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[496] ),
        .I2(\f_permutation_l_/out_reg_n_0_[71] ),
        .I3(\out[1500]_i_3_n_0 ),
        .I4(\out[639]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [447]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[448]_i_1 
       (.I0(\out[1570]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[886] ),
        .I2(\out[448]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[72] ),
        .I4(\out[1501]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [448]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[448]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[497] ),
        .I1(\f_permutation_l_/round_in [1392]),
        .I2(\out[1564]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1521]),
        .I4(\out[1564]_i_9_n_0 ),
        .O(\out[448]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[449]_i_1 
       (.I0(\out[1571]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[887] ),
        .I2(\out[449]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[73] ),
        .I4(\out[1502]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [449]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[449]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[498] ),
        .I1(\f_permutation_l_/round_in [1393]),
        .I2(\out[1565]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1522]),
        .I4(\out[1565]_i_9_n_0 ),
        .O(\out[449]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[44]_i_1 
       (.I0(\out[1558]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[234] ),
        .I2(\out[300]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1077]),
        .I4(\out[1482]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[450]_i_1 
       (.I0(\out[1572]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[888] ),
        .I2(\out[450]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[74] ),
        .I4(\out[1503]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [450]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[450]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[499] ),
        .I1(\f_permutation_l_/round_in [1394]),
        .I2(\out[1566]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1523]),
        .I4(\out[1566]_i_9_n_0 ),
        .O(\out[450]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[451]_i_1 
       (.I0(\out[1573]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[889] ),
        .I2(\out[451]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[75] ),
        .I4(\out[1504]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [451]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[451]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[500] ),
        .I1(\f_permutation_l_/round_in [1395]),
        .I2(\out[1567]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1524]),
        .I4(\out[1567]_i_10_n_0 ),
        .O(\out[451]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[452]_i_1 
       (.I0(\out[1574]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[890] ),
        .I2(\out[452]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[76] ),
        .I4(\out[1505]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [452]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[452]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[501] ),
        .I1(\f_permutation_l_/round_in [1396]),
        .I2(\out[1568]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1525]),
        .I4(\out[1568]_i_9_n_0 ),
        .O(\out[452]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[453]_i_1 
       (.I0(\out[1575]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[891] ),
        .I2(\out[453]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[77] ),
        .I4(\out[1506]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [453]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[453]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[502] ),
        .I1(\f_permutation_l_/round_in [1397]),
        .I2(\out[1569]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1526]),
        .I4(\out[1569]_i_9_n_0 ),
        .O(\out[453]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[454]_i_1 
       (.I0(\out[1576]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[892] ),
        .I2(\out[454]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[78] ),
        .I4(\out[1507]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [454]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[454]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[503] ),
        .I1(\f_permutation_l_/round_in [1398]),
        .I2(\out[1570]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1527]),
        .I4(\out[1570]_i_9_n_0 ),
        .O(\out[454]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[455]_i_1 
       (.I0(\out[1577]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[893] ),
        .I2(\out[455]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[79] ),
        .I4(\out[1508]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [455]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[455]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[504] ),
        .I1(\f_permutation_l_/round_in [1399]),
        .I2(\out[1571]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1528]),
        .I4(\out[1571]_i_9_n_0 ),
        .O(\out[455]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[456]_i_1 
       (.I0(\out[1578]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[894] ),
        .I2(\out[456]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[80] ),
        .I4(\out[1509]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [456]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[456]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[505] ),
        .I1(\f_permutation_l_/round_in [1400]),
        .I2(\out[1572]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1529]),
        .I4(\out[1572]_i_9_n_0 ),
        .O(\out[456]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[457]_i_1 
       (.I0(\out[1579]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[895] ),
        .I2(\out[457]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[81] ),
        .I4(\out[1510]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [457]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[457]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[506] ),
        .I1(\f_permutation_l_/round_in [1401]),
        .I2(\out[1573]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1530]),
        .I4(\out[1573]_i_9_n_0 ),
        .O(\out[457]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[458]_i_1 
       (.I0(\out[1580]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[832] ),
        .I2(\out[458]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[82] ),
        .I4(\out[1511]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [458]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[458]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[507] ),
        .I1(\f_permutation_l_/round_in [1402]),
        .I2(\out[1574]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1531]),
        .I4(\out[1574]_i_9_n_0 ),
        .O(\out[458]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[459]_i_1 
       (.I0(\out[1581]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[833] ),
        .I2(\out[459]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[83] ),
        .I4(\out[1512]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [459]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[459]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[508] ),
        .I1(\f_permutation_l_/round_in [1403]),
        .I2(\out[1575]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1532]),
        .I4(\out[1575]_i_9_n_0 ),
        .O(\out[459]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[45]_i_1 
       (.I0(\out[1559]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[235] ),
        .I2(\out[301]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1078]),
        .I4(\out[1483]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[460]_i_1 
       (.I0(\out[1582]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[834] ),
        .I2(\out[460]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[84] ),
        .I4(\out[1513]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [460]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[460]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[509] ),
        .I1(\f_permutation_l_/round_in [1404]),
        .I2(\out[1576]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1533]),
        .I4(\out[1576]_i_9_n_0 ),
        .O(\out[460]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[461]_i_1 
       (.I0(\out[1583]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[835] ),
        .I2(\out[461]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[85] ),
        .I4(\out[1514]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [461]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[461]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[510] ),
        .I1(\f_permutation_l_/round_in [1405]),
        .I2(\out[1577]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1534]),
        .I4(\out[1577]_i_9_n_0 ),
        .O(\out[461]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[462]_i_1 
       (.I0(\out[1584]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[836] ),
        .I2(\out[462]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[86] ),
        .I4(\out[1515]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [462]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[462]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[511] ),
        .I1(\f_permutation_l_/round_in [1406]),
        .I2(\out[1578]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[462]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[463]_i_1 
       (.I0(\out[1585]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[837] ),
        .I2(\out[463]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[87] ),
        .I4(\out[1516]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [463]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[463]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[448] ),
        .I1(\f_permutation_l_/round_in [1407]),
        .I2(\out[1579]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[463]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[464]_i_1 
       (.I0(\out[1586]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[838] ),
        .I2(\out[464]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[88] ),
        .I4(\out[1517]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [464]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[464]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[449] ),
        .I1(\f_permutation_l_/round_in [1344]),
        .I2(\out[1580]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[464]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[465]_i_1 
       (.I0(\out[1587]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[839] ),
        .I2(\out[465]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[89] ),
        .I4(\out[1518]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [465]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[465]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[450] ),
        .I1(\f_permutation_l_/round_in [1345]),
        .I2(\out[1581]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[465]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[466]_i_1 
       (.I0(\out[1588]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[840] ),
        .I2(\out[466]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[90] ),
        .I4(\out[1519]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [466]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[466]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[451] ),
        .I1(\f_permutation_l_/round_in [1346]),
        .I2(\out[1582]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[466]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[467]_i_1 
       (.I0(\out[1589]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[841] ),
        .I2(\out[467]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[91] ),
        .I4(\out[1520]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [467]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[467]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[452] ),
        .I1(\f_permutation_l_/round_in [1347]),
        .I2(\out[1583]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[467]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[468]_i_1 
       (.I0(\out[1590]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[842] ),
        .I2(\out[468]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[92] ),
        .I4(\out[1521]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [468]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[468]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[453] ),
        .I1(\f_permutation_l_/round_in [1348]),
        .I2(\out[1584]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[468]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[469]_i_1 
       (.I0(\out[1591]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[843] ),
        .I2(\out[469]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[93] ),
        .I4(\out[1522]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [469]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[469]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[454] ),
        .I1(\f_permutation_l_/round_in [1349]),
        .I2(\out[1585]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[469]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[46]_i_1 
       (.I0(\out[1560]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[236] ),
        .I2(\out[302]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1079]),
        .I4(\out[1484]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[470]_i_1 
       (.I0(\out[1592]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[844] ),
        .I2(\out[470]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[94] ),
        .I4(\out[1523]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [470]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[470]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[455] ),
        .I1(\f_permutation_l_/round_in [1350]),
        .I2(\out[1586]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[470]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[471]_i_1 
       (.I0(\out[1593]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[845] ),
        .I2(\out[471]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[95] ),
        .I4(\out[1524]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [471]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[471]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[456] ),
        .I1(\f_permutation_l_/round_in [1351]),
        .I2(\out[1587]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[471]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[472]_i_1 
       (.I0(\out[1594]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[846] ),
        .I2(\out[472]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[96] ),
        .I4(\out[1525]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [472]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[472]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[457] ),
        .I1(\f_permutation_l_/round_in [1352]),
        .I2(\out[1588]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[472]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[473]_i_1 
       (.I0(\out[1595]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[847] ),
        .I2(\out[473]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[97] ),
        .I4(\out[1526]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [473]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[473]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[458] ),
        .I1(\f_permutation_l_/round_in [1353]),
        .I2(\out[1589]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[473]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[474]_i_1 
       (.I0(\out[1596]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[848] ),
        .I2(\out[474]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[98] ),
        .I4(\out[1527]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [474]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[474]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[459] ),
        .I1(\f_permutation_l_/round_in [1354]),
        .I2(\out[1590]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[474]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[475]_i_1 
       (.I0(\out[1597]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[849] ),
        .I2(\out[475]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[99] ),
        .I4(\out[1528]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [475]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[475]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[460] ),
        .I1(\f_permutation_l_/round_in [1355]),
        .I2(\out[1591]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[475]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[476]_i_1 
       (.I0(\out[1598]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[850] ),
        .I2(\out[476]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[100] ),
        .I4(\out[1529]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [476]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[476]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[461] ),
        .I1(\f_permutation_l_/round_in [1356]),
        .I2(\out[1592]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[476]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[477]_i_1 
       (.I0(\out[1343]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[851] ),
        .I2(\out[477]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[101] ),
        .I4(\out[1530]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [477]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[477]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[462] ),
        .I1(\f_permutation_l_/round_in [1357]),
        .I2(\out[1593]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[477]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[478]_i_1 
       (.I0(\out[1280]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[852] ),
        .I2(\out[478]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[102] ),
        .I4(\out[1531]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [478]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[478]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[463] ),
        .I1(\f_permutation_l_/round_in [1358]),
        .I2(\out[1594]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[478]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[479]_i_1 
       (.I0(\out[1281]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[853] ),
        .I2(\out[479]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[103] ),
        .I4(\out[1532]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [479]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[479]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[464] ),
        .I1(\f_permutation_l_/round_in [1359]),
        .I2(\out[1595]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[479]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[47]_i_1 
       (.I0(\out[1561]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[237] ),
        .I2(\out[303]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1080]),
        .I4(\out[1485]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[480]_i_1 
       (.I0(\out[1538]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[854] ),
        .I2(\out[480]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[104] ),
        .I4(\out[1533]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [480]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[480]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[465] ),
        .I1(\f_permutation_l_/round_in [1360]),
        .I2(\out[1596]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[480]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[481]_i_1 
       (.I0(\out[1539]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[855] ),
        .I2(\out[481]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[105] ),
        .I4(\out[1534]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [481]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[481]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[466] ),
        .I1(\f_permutation_l_/round_in [1361]),
        .I2(\out[1597]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[481]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[482]_i_1 
       (.I0(\out[1540]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[856] ),
        .I2(\out[482]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[106] ),
        .I4(\out[1535]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [482]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[482]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[467] ),
        .I1(\f_permutation_l_/round_in [1362]),
        .I2(\out[1598]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[482]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[483]_i_1 
       (.I0(\out[1541]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[857] ),
        .I2(\out[483]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[107] ),
        .I4(\out[1472]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [483]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[483]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[468] ),
        .I1(\f_permutation_l_/round_in [1363]),
        .I2(\out[1599]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[483]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[484]_i_1 
       (.I0(\out[1542]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[858] ),
        .I2(\out[484]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[108] ),
        .I4(\out[1473]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [484]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[484]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[469] ),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1493]),
        .I4(\out[1536]_i_14_n_0 ),
        .O(\out[484]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[485]_i_1 
       (.I0(\out[1287]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[859] ),
        .I2(\out[485]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[109] ),
        .I4(\out[1474]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [485]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[485]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[470] ),
        .I1(\f_permutation_l_/round_in [1365]),
        .I2(\out[1537]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1494]),
        .I4(\out[1537]_i_10_n_0 ),
        .O(\out[485]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[486]_i_1 
       (.I0(\out[1544]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[860] ),
        .I2(\out[486]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[110] ),
        .I4(\out[1475]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [486]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[486]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[471] ),
        .I1(\f_permutation_l_/round_in [1366]),
        .I2(\out[1538]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1495]),
        .I4(\out[1538]_i_9_n_0 ),
        .O(\out[486]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[487]_i_1 
       (.I0(\out[1545]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[861] ),
        .I2(\out[487]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[111] ),
        .I4(\out[1476]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [487]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[487]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[472] ),
        .I1(\out[1539]_i_12_n_0 ),
        .I2(\f_permutation_l_/round_in [1367]),
        .I3(\f_permutation_l_/round_in [1496]),
        .I4(\out[1539]_i_14_n_0 ),
        .O(\out[487]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[488]_i_1 
       (.I0(\out[1546]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[862] ),
        .I2(\out[488]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[112] ),
        .I4(\out[1477]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [488]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[488]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[473] ),
        .I1(\f_permutation_l_/round_in [1368]),
        .I2(\out[1540]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1497]),
        .I4(\out[1540]_i_9_n_0 ),
        .O(\out[488]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[489]_i_1 
       (.I0(\out[1547]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[863] ),
        .I2(\out[489]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[113] ),
        .I4(\out[1478]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [489]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[489]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[474] ),
        .I1(\f_permutation_l_/round_in [1369]),
        .I2(\out[1541]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1498]),
        .I4(\out[1541]_i_9_n_0 ),
        .O(\out[489]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[48]_i_1 
       (.I0(\out[1562]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[238] ),
        .I2(\out[304]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1081]),
        .I4(\out[1486]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[490]_i_1 
       (.I0(\out[1548]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[864] ),
        .I2(\out[490]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[114] ),
        .I4(\out[1479]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [490]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[490]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[475] ),
        .I1(\f_permutation_l_/round_in [1370]),
        .I2(\out[1542]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1499]),
        .I4(\out[1542]_i_11_n_0 ),
        .O(\out[490]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[491]_i_1 
       (.I0(\out[1549]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[865] ),
        .I2(\out[491]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[115] ),
        .I4(\out[1480]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [491]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[491]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[476] ),
        .I1(\f_permutation_l_/round_in [1371]),
        .I2(\out[1543]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1500]),
        .I4(\out[1543]_i_11_n_0 ),
        .O(\out[491]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[492]_i_1 
       (.I0(\out[1550]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[866] ),
        .I2(\out[492]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[116] ),
        .I4(\out[1481]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [492]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[492]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[477] ),
        .I1(\f_permutation_l_/round_in [1372]),
        .I2(\out[1544]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1501]),
        .I4(\out[1544]_i_9_n_0 ),
        .O(\out[492]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[493]_i_1 
       (.I0(\out[1295]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[867] ),
        .I2(\out[493]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[117] ),
        .I4(\out[1482]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [493]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[493]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[478] ),
        .I1(\f_permutation_l_/round_in [1373]),
        .I2(\out[1545]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1502]),
        .I4(\out[1545]_i_9_n_0 ),
        .O(\out[493]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[494]_i_1 
       (.I0(\out[1552]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[868] ),
        .I2(\out[494]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[118] ),
        .I4(\out[1483]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [494]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[494]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[479] ),
        .I1(\f_permutation_l_/round_in [1374]),
        .I2(\out[1546]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1503]),
        .I4(\out[1546]_i_9_n_0 ),
        .O(\out[494]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[495]_i_1 
       (.I0(\out[1553]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[869] ),
        .I2(\out[495]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[119] ),
        .I4(\out[1484]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [495]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[495]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[480] ),
        .I1(\f_permutation_l_/round_in [1375]),
        .I2(\out[1547]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1504]),
        .I4(\out[1547]_i_9_n_0 ),
        .O(\out[495]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[496]_i_1 
       (.I0(\out[1554]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[870] ),
        .I2(\out[496]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[120] ),
        .I4(\out[1485]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [496]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[496]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[481] ),
        .I1(\f_permutation_l_/round_in [1376]),
        .I2(\out[1548]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1505]),
        .I4(\out[1548]_i_9_n_0 ),
        .O(\out[496]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[497]_i_1 
       (.I0(\out[1555]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[871] ),
        .I2(\out[497]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[121] ),
        .I4(\out[1486]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [497]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[497]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[482] ),
        .I1(\f_permutation_l_/round_in [1377]),
        .I2(\out[1549]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1506]),
        .I4(\out[1549]_i_9_n_0 ),
        .O(\out[497]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[498]_i_1 
       (.I0(\out[1556]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[872] ),
        .I2(\out[498]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[122] ),
        .I4(\out[1487]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [498]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[498]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[483] ),
        .I1(\f_permutation_l_/round_in [1378]),
        .I2(\out[1550]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1507]),
        .I4(\out[1550]_i_9_n_0 ),
        .O(\out[498]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[499]_i_1 
       (.I0(\out[1557]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[873] ),
        .I2(\out[499]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[123] ),
        .I4(\out[1488]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [499]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[499]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[484] ),
        .I1(\f_permutation_l_/round_in [1379]),
        .I2(\out[1551]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1508]),
        .I4(\out[1551]_i_10_n_0 ),
        .O(\out[499]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[49]_i_1 
       (.I0(\out[1563]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[239] ),
        .I2(\out[305]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1082]),
        .I4(\out[1487]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[4]_i_1 
       (.I0(\out[1582]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[194] ),
        .I2(\out[260]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1037]),
        .I4(\out[1506]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[500]_i_1 
       (.I0(\out[1558]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[874] ),
        .I2(\out[500]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[124] ),
        .I4(\out[1489]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [500]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[500]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[485] ),
        .I1(\f_permutation_l_/round_in [1380]),
        .I2(\out[1552]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1509]),
        .I4(\out[1552]_i_9_n_0 ),
        .O(\out[500]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[501]_i_1 
       (.I0(\out[1559]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[875] ),
        .I2(\out[501]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[125] ),
        .I4(\out[1490]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [501]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[501]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[486] ),
        .I1(\f_permutation_l_/round_in [1381]),
        .I2(\out[1553]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1510]),
        .I4(\out[1553]_i_9_n_0 ),
        .O(\out[501]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[502]_i_1 
       (.I0(\out[1560]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[876] ),
        .I2(\out[502]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[126] ),
        .I4(\out[1491]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [502]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[502]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[487] ),
        .I1(\f_permutation_l_/round_in [1382]),
        .I2(\out[1554]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1511]),
        .I4(\out[1554]_i_9_n_0 ),
        .O(\out[502]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[503]_i_1 
       (.I0(\out[1561]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[877] ),
        .I2(\out[503]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[127] ),
        .I4(\out[1492]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [503]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[503]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[488] ),
        .I1(\f_permutation_l_/round_in [1383]),
        .I2(\out[1555]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1512]),
        .I4(\out[1555]_i_9_n_0 ),
        .O(\out[503]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[504]_i_1 
       (.I0(\out[1562]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[878] ),
        .I2(\out[504]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[64] ),
        .I4(\out[1493]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [504]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[504]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[489] ),
        .I1(\f_permutation_l_/round_in [1384]),
        .I2(\out[1556]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1513]),
        .I4(\out[1556]_i_10_n_0 ),
        .O(\out[504]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[505]_i_1 
       (.I0(\out[1563]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[879] ),
        .I2(\out[505]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[65] ),
        .I4(\out[1494]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [505]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[505]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[490] ),
        .I1(\f_permutation_l_/round_in [1385]),
        .I2(\out[1557]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1514]),
        .I4(\out[1557]_i_9_n_0 ),
        .O(\out[505]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[506]_i_1 
       (.I0(\out[1564]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[880] ),
        .I2(\out[506]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[66] ),
        .I4(\out[1495]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [506]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[506]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[491] ),
        .I1(\f_permutation_l_/round_in [1386]),
        .I2(\out[1558]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1515]),
        .I4(\out[1558]_i_9_n_0 ),
        .O(\out[506]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[507]_i_1 
       (.I0(\out[1565]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[881] ),
        .I2(\out[507]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[67] ),
        .I4(\out[1496]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [507]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[507]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[492] ),
        .I1(\f_permutation_l_/round_in [1387]),
        .I2(\out[1559]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1516]),
        .I4(\out[1559]_i_9_n_0 ),
        .O(\out[507]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[508]_i_1 
       (.I0(\out[1566]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[882] ),
        .I2(\out[508]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[68] ),
        .I4(\out[1497]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [508]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[508]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[493] ),
        .I1(\f_permutation_l_/round_in [1388]),
        .I2(\out[1560]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1517]),
        .I4(\out[1560]_i_9_n_0 ),
        .O(\out[508]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[509]_i_1 
       (.I0(\out[1311]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[883] ),
        .I2(\out[509]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[69] ),
        .I4(\out[1498]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [509]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[509]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[494] ),
        .I1(\f_permutation_l_/round_in [1389]),
        .I2(\out[1561]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1518]),
        .I4(\out[1561]_i_9_n_0 ),
        .O(\out[509]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[50]_i_1 
       (.I0(\out[1564]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[240] ),
        .I2(\out[306]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1083]),
        .I4(\out[1488]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[510]_i_1 
       (.I0(\out[1568]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[884] ),
        .I2(\out[510]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[70] ),
        .I4(\out[1499]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [510]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[510]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[495] ),
        .I1(\f_permutation_l_/round_in [1390]),
        .I2(\out[1562]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1519]),
        .I4(\out[1562]_i_9_n_0 ),
        .O(\out[510]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[511]_i_1 
       (.I0(\out[1569]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[885] ),
        .I2(\out[511]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[71] ),
        .I4(\out[1500]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [511]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[511]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[496] ),
        .I1(\f_permutation_l_/round_in [1391]),
        .I2(\out[1563]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1520]),
        .I4(\out[1563]_i_9_n_0 ),
        .O(\out[511]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[512]_i_1 
       (.I0(\out[512]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[886] ),
        .I2(\out[1570]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[497] ),
        .I4(\out[1564]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [512]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[512]_i_2 
       (.I0(\f_permutation_l_/round_in [1244]),
        .I1(\f_permutation_l_/round_in [1499]),
        .I2(\out[1542]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1308]),
        .I4(\out[1564]_i_15_n_0 ),
        .O(\out[512]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[513]_i_1 
       (.I0(\out[513]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[887] ),
        .I2(\out[1571]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[498] ),
        .I4(\out[1565]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [513]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[513]_i_2 
       (.I0(\f_permutation_l_/round_in [1245]),
        .I1(\f_permutation_l_/round_in [1500]),
        .I2(\out[1543]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1309]),
        .I4(\out[1565]_i_15_n_0 ),
        .O(\out[513]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[514]_i_1 
       (.I0(\out[514]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[888] ),
        .I2(\out[1572]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[499] ),
        .I4(\out[1566]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [514]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[514]_i_2 
       (.I0(\f_permutation_l_/round_in [1246]),
        .I1(\f_permutation_l_/round_in [1501]),
        .I2(\out[1544]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1310]),
        .I4(\out[1566]_i_14_n_0 ),
        .O(\out[514]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[515]_i_1 
       (.I0(\out[515]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[889] ),
        .I2(\out[1573]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[500] ),
        .I4(\out[1567]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [515]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[515]_i_2 
       (.I0(\f_permutation_l_/round_in [1247]),
        .I1(\f_permutation_l_/round_in [1502]),
        .I2(\out[1545]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1311]),
        .I4(\out[1567]_i_16_n_0 ),
        .O(\out[515]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[516]_i_1 
       (.I0(\out[516]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[890] ),
        .I2(\out[1574]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[501] ),
        .I4(\out[1568]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [516]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[516]_i_2 
       (.I0(\f_permutation_l_/round_in [1248]),
        .I1(\f_permutation_l_/round_in [1503]),
        .I2(\out[1546]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1312]),
        .I4(\out[1568]_i_15_n_0 ),
        .O(\out[516]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[517]_i_1 
       (.I0(\out[517]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[891] ),
        .I2(\out[1575]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[502] ),
        .I4(\out[1569]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [517]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[517]_i_2 
       (.I0(\f_permutation_l_/round_in [1249]),
        .I1(\f_permutation_l_/round_in [1504]),
        .I2(\out[1547]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1313]),
        .I4(\out[1569]_i_15_n_0 ),
        .O(\out[517]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[518]_i_1 
       (.I0(\out[518]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[892] ),
        .I2(\out[1576]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[503] ),
        .I4(\out[1570]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [518]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[518]_i_2 
       (.I0(\f_permutation_l_/round_in [1250]),
        .I1(\f_permutation_l_/round_in [1505]),
        .I2(\out[1548]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1314]),
        .I4(\out[1570]_i_15_n_0 ),
        .O(\out[518]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[519]_i_1 
       (.I0(\out[519]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[893] ),
        .I2(\out[1577]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[504] ),
        .I4(\out[1571]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [519]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[519]_i_2 
       (.I0(\f_permutation_l_/round_in [1251]),
        .I1(\f_permutation_l_/round_in [1506]),
        .I2(\out[1549]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1315]),
        .I4(\out[1571]_i_14_n_0 ),
        .O(\out[519]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[51]_i_1 
       (.I0(\out[1565]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[241] ),
        .I2(\out[307]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1084]),
        .I4(\out[1489]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[520]_i_1 
       (.I0(\out[520]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[894] ),
        .I2(\out[1578]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[505] ),
        .I4(\out[1572]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [520]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[520]_i_2 
       (.I0(\f_permutation_l_/round_in [1252]),
        .I1(\f_permutation_l_/round_in [1507]),
        .I2(\out[1550]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1316]),
        .I4(\out[1572]_i_15_n_0 ),
        .O(\out[520]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[521]_i_1 
       (.I0(\out[521]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[895] ),
        .I2(\out[1579]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[506] ),
        .I4(\out[1573]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [521]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[521]_i_2 
       (.I0(\f_permutation_l_/round_in [1253]),
        .I1(\f_permutation_l_/round_in [1508]),
        .I2(\out[1551]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1317]),
        .I4(\out[1573]_i_15_n_0 ),
        .O(\out[521]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[522]_i_1 
       (.I0(\out[522]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[832] ),
        .I2(\out[1580]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[507] ),
        .I4(\out[1574]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [522]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[522]_i_2 
       (.I0(\f_permutation_l_/round_in [1254]),
        .I1(\f_permutation_l_/round_in [1509]),
        .I2(\out[1552]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1318]),
        .I4(\out[1574]_i_15_n_0 ),
        .O(\out[522]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[523]_i_1 
       (.I0(\out[523]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[833] ),
        .I2(\out[1581]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[508] ),
        .I4(\out[1575]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [523]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[523]_i_2 
       (.I0(\f_permutation_l_/round_in [1255]),
        .I1(\f_permutation_l_/round_in [1510]),
        .I2(\out[1553]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1319]),
        .I4(\out[1575]_i_15_n_0 ),
        .O(\out[523]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[524]_i_1 
       (.I0(\out[524]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[834] ),
        .I2(\out[1582]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[509] ),
        .I4(\out[1576]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [524]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[524]_i_2 
       (.I0(\f_permutation_l_/round_in [1256]),
        .I1(\f_permutation_l_/round_in [1511]),
        .I2(\out[1554]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1320]),
        .I4(\out[1576]_i_15_n_0 ),
        .O(\out[524]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[525]_i_1 
       (.I0(\out[525]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[835] ),
        .I2(\out[1583]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[510] ),
        .I4(\out[1577]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [525]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[525]_i_2 
       (.I0(\f_permutation_l_/round_in [1257]),
        .I1(\f_permutation_l_/round_in [1512]),
        .I2(\out[1555]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1321]),
        .I4(\out[1577]_i_15_n_0 ),
        .O(\out[525]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[526]_i_1 
       (.I0(\out[526]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[836] ),
        .I2(\out[1584]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[511] ),
        .I4(\out[1578]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [526]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[526]_i_2 
       (.I0(\f_permutation_l_/round_in [1258]),
        .I1(\f_permutation_l_/round_in [1513]),
        .I2(\out[1556]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1322]),
        .I4(\out[1578]_i_14_n_0 ),
        .O(\out[526]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[527]_i_1 
       (.I0(\out[527]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[837] ),
        .I2(\out[1585]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[448] ),
        .I4(\out[1579]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [527]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[527]_i_2 
       (.I0(\f_permutation_l_/round_in [1259]),
        .I1(\f_permutation_l_/round_in [1514]),
        .I2(\out[1557]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1323]),
        .I4(\out[1579]_i_15_n_0 ),
        .O(\out[527]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[528]_i_1 
       (.I0(\out[528]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[838] ),
        .I2(\out[1586]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[449] ),
        .I4(\out[1580]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [528]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[528]_i_2 
       (.I0(\f_permutation_l_/round_in [1260]),
        .I1(\f_permutation_l_/round_in [1515]),
        .I2(\out[1558]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1324]),
        .I4(\out[1580]_i_14_n_0 ),
        .O(\out[528]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[529]_i_1 
       (.I0(\out[529]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[839] ),
        .I2(\out[1587]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[450] ),
        .I4(\out[1581]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [529]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[529]_i_2 
       (.I0(\f_permutation_l_/round_in [1261]),
        .I1(\f_permutation_l_/round_in [1516]),
        .I2(\out[1559]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1325]),
        .I4(\out[1581]_i_14_n_0 ),
        .O(\out[529]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[52]_i_1 
       (.I0(\out[1566]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[242] ),
        .I2(\out[308]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1085]),
        .I4(\out[1490]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[530]_i_1 
       (.I0(\out[530]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[840] ),
        .I2(\out[1588]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[451] ),
        .I4(\out[1582]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [530]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[530]_i_2 
       (.I0(\f_permutation_l_/round_in [1262]),
        .I1(\f_permutation_l_/round_in [1517]),
        .I2(\out[1560]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1326]),
        .I4(\out[1582]_i_14_n_0 ),
        .O(\out[530]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[531]_i_1 
       (.I0(\out[531]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[841] ),
        .I2(\out[1589]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[452] ),
        .I4(\out[1583]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [531]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[531]_i_2 
       (.I0(\f_permutation_l_/round_in [1263]),
        .I1(\f_permutation_l_/round_in [1518]),
        .I2(\out[1561]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1327]),
        .I4(\out[1583]_i_14_n_0 ),
        .O(\out[531]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[532]_i_1 
       (.I0(\out[532]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[842] ),
        .I2(\out[1590]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[453] ),
        .I4(\out[1584]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [532]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[532]_i_2 
       (.I0(\f_permutation_l_/round_in [1264]),
        .I1(\f_permutation_l_/round_in [1519]),
        .I2(\out[1562]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1328]),
        .I4(\out[1584]_i_14_n_0 ),
        .O(\out[532]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[533]_i_1 
       (.I0(\out[533]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[843] ),
        .I2(\out[1591]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[454] ),
        .I4(\out[1585]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [533]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[533]_i_2 
       (.I0(\f_permutation_l_/round_in [1265]),
        .I1(\f_permutation_l_/round_in [1520]),
        .I2(\out[1563]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1329]),
        .I4(\out[1585]_i_14_n_0 ),
        .O(\out[533]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[534]_i_1 
       (.I0(\out[534]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[844] ),
        .I2(\out[1592]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[455] ),
        .I4(\out[1586]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [534]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[534]_i_2 
       (.I0(\f_permutation_l_/round_in [1266]),
        .I1(\f_permutation_l_/round_in [1521]),
        .I2(\out[1564]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1330]),
        .I4(\out[1586]_i_14_n_0 ),
        .O(\out[534]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[535]_i_1 
       (.I0(\out[535]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[845] ),
        .I2(\out[1593]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[456] ),
        .I4(\out[1587]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [535]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[535]_i_2 
       (.I0(\f_permutation_l_/round_in [1267]),
        .I1(\f_permutation_l_/round_in [1522]),
        .I2(\out[1565]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1331]),
        .I4(\out[1587]_i_13_n_0 ),
        .O(\out[535]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[536]_i_1 
       (.I0(\out[536]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[846] ),
        .I2(\out[1594]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[457] ),
        .I4(\out[1588]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [536]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[536]_i_2 
       (.I0(\f_permutation_l_/round_in [1268]),
        .I1(\f_permutation_l_/round_in [1523]),
        .I2(\out[1566]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1332]),
        .I4(\out[1588]_i_14_n_0 ),
        .O(\out[536]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[537]_i_1 
       (.I0(\out[537]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[847] ),
        .I2(\out[1595]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[458] ),
        .I4(\out[1589]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [537]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[537]_i_2 
       (.I0(\f_permutation_l_/round_in [1269]),
        .I1(\f_permutation_l_/round_in [1524]),
        .I2(\out[1567]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1333]),
        .I4(\out[1589]_i_14_n_0 ),
        .O(\out[537]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[538]_i_1 
       (.I0(\out[538]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[848] ),
        .I2(\out[1596]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[459] ),
        .I4(\out[1590]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [538]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[538]_i_2 
       (.I0(\f_permutation_l_/round_in [1270]),
        .I1(\f_permutation_l_/round_in [1525]),
        .I2(\out[1568]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1334]),
        .I4(\out[1590]_i_14_n_0 ),
        .O(\out[538]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[539]_i_1 
       (.I0(\out[539]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[849] ),
        .I2(\out[1597]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[460] ),
        .I4(\out[1591]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [539]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[539]_i_2 
       (.I0(\f_permutation_l_/round_in [1271]),
        .I1(\f_permutation_l_/round_in [1526]),
        .I2(\out[1569]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1335]),
        .I4(\out[1591]_i_14_n_0 ),
        .O(\out[539]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[53]_i_1 
       (.I0(\out[1311]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[243] ),
        .I2(\out[309]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1086]),
        .I4(\out[1491]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[540]_i_1 
       (.I0(\out[540]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[850] ),
        .I2(\out[1598]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[461] ),
        .I4(\out[1592]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [540]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[540]_i_2 
       (.I0(\f_permutation_l_/round_in [1272]),
        .I1(\f_permutation_l_/round_in [1527]),
        .I2(\out[1570]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1336]),
        .I4(\out[1592]_i_14_n_0 ),
        .O(\out[540]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[541]_i_1 
       (.I0(\out[541]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[851] ),
        .I2(\out[1343]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[462] ),
        .I4(\out[1593]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [541]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[541]_i_2 
       (.I0(\f_permutation_l_/round_in [1273]),
        .I1(\f_permutation_l_/round_in [1528]),
        .I2(\out[1571]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1337]),
        .I4(\out[1593]_i_14_n_0 ),
        .O(\out[541]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[542]_i_1 
       (.I0(\out[542]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[852] ),
        .I2(\out[1280]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[463] ),
        .I4(\out[1594]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [542]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[542]_i_2 
       (.I0(\f_permutation_l_/round_in [1274]),
        .I1(\f_permutation_l_/round_in [1529]),
        .I2(\out[1572]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1338]),
        .I4(\out[1594]_i_14_n_0 ),
        .O(\out[542]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[543]_i_1 
       (.I0(\out[543]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[853] ),
        .I2(\out[1281]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[464] ),
        .I4(\out[1595]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [543]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[543]_i_2 
       (.I0(\f_permutation_l_/round_in [1275]),
        .I1(\f_permutation_l_/round_in [1530]),
        .I2(\out[1573]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1339]),
        .I4(\out[1595]_i_14_n_0 ),
        .O(\out[543]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[544]_i_1 
       (.I0(\out[544]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[854] ),
        .I2(\out[1538]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[465] ),
        .I4(\out[1596]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [544]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[544]_i_2 
       (.I0(\f_permutation_l_/round_in [1276]),
        .I1(\f_permutation_l_/round_in [1531]),
        .I2(\out[1574]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1340]),
        .I4(\out[1596]_i_14_n_0 ),
        .O(\out[544]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[545]_i_1 
       (.I0(\out[545]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[855] ),
        .I2(\out[1539]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[466] ),
        .I4(\out[1597]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [545]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[545]_i_2 
       (.I0(\f_permutation_l_/round_in [1277]),
        .I1(\f_permutation_l_/round_in [1532]),
        .I2(\out[1575]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1341]),
        .I4(\out[1597]_i_14_n_0 ),
        .O(\out[545]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[546]_i_1 
       (.I0(\out[546]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[856] ),
        .I2(\out[1540]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[467] ),
        .I4(\out[1598]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [546]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[546]_i_2 
       (.I0(\f_permutation_l_/round_in [1278]),
        .I1(\f_permutation_l_/round_in [1533]),
        .I2(\out[1576]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1342]),
        .I4(\out[1598]_i_14_n_0 ),
        .O(\out[546]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[547]_i_1 
       (.I0(\out[547]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[857] ),
        .I2(\out[1541]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[468] ),
        .I4(\out[1599]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [547]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[547]_i_2 
       (.I0(\f_permutation_l_/round_in [1279]),
        .I1(\f_permutation_l_/round_in [1534]),
        .I2(\out[1577]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1343]),
        .I4(\out[1599]_i_14_n_0 ),
        .O(\out[547]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[548]_i_1 
       (.I0(\out[548]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[858] ),
        .I2(\out[1542]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[469] ),
        .I4(\out[1472]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [548]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[548]_i_2 
       (.I0(\f_permutation_l_/round_in [1216]),
        .I1(\f_permutation_l_/round_in [1280]),
        .I2(\out[1536]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[548]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[549]_i_1 
       (.I0(\out[549]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[859] ),
        .I2(\out[1287]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[470] ),
        .I4(\out[1537]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [549]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[549]_i_2 
       (.I0(\f_permutation_l_/round_in [1217]),
        .I1(\f_permutation_l_/round_in [1281]),
        .I2(\out[1537]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[549]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[54]_i_1 
       (.I0(\out[1568]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[244] ),
        .I2(\out[310]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1087]),
        .I4(\out[1492]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[550]_i_1 
       (.I0(\out[550]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[860] ),
        .I2(\out[1544]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[471] ),
        .I4(\out[1538]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [550]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[550]_i_2 
       (.I0(\f_permutation_l_/round_in [1218]),
        .I1(\f_permutation_l_/round_in [1282]),
        .I2(\out[1538]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[550]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[551]_i_1 
       (.I0(\out[551]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[861] ),
        .I2(\out[1545]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[472] ),
        .I4(\out[1045]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [551]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[551]_i_2 
       (.I0(\f_permutation_l_/round_in [1219]),
        .I1(\f_permutation_l_/round_in [1283]),
        .I2(\out[1539]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[551]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[552]_i_1 
       (.I0(\out[552]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[862] ),
        .I2(\out[1546]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[473] ),
        .I4(\out[1540]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [552]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[552]_i_2 
       (.I0(\f_permutation_l_/round_in [1220]),
        .I1(\f_permutation_l_/round_in [1284]),
        .I2(\out[1540]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[552]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[553]_i_1 
       (.I0(\out[553]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[863] ),
        .I2(\out[1547]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[474] ),
        .I4(\out[1541]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [553]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[553]_i_2 
       (.I0(\f_permutation_l_/round_in [1221]),
        .I1(\f_permutation_l_/round_in [1285]),
        .I2(\out[1541]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[553]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[554]_i_1 
       (.I0(\out[554]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[864] ),
        .I2(\out[1548]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[475] ),
        .I4(\out[1542]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [554]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[554]_i_2 
       (.I0(\f_permutation_l_/round_in [1222]),
        .I1(\f_permutation_l_/round_in [1286]),
        .I2(\out[1542]_i_16_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[554]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[555]_i_1 
       (.I0(\out[555]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[865] ),
        .I2(\out[1549]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[476] ),
        .I4(\out[1543]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [555]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[555]_i_2 
       (.I0(\f_permutation_l_/round_in [1223]),
        .I1(\f_permutation_l_/round_in [1287]),
        .I2(\out[1543]_i_17_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[555]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[556]_i_1 
       (.I0(\out[556]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[866] ),
        .I2(\out[1550]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[477] ),
        .I4(\out[1544]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [556]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[556]_i_2 
       (.I0(\f_permutation_l_/round_in [1224]),
        .I1(\f_permutation_l_/round_in [1288]),
        .I2(\out[1544]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[556]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[557]_i_1 
       (.I0(\out[557]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[867] ),
        .I2(\out[1295]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[478] ),
        .I4(\out[1545]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [557]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[557]_i_2 
       (.I0(\f_permutation_l_/round_in [1225]),
        .I1(\f_permutation_l_/round_in [1289]),
        .I2(\out[1545]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[557]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[558]_i_1 
       (.I0(\out[558]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[868] ),
        .I2(\out[1552]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[479] ),
        .I4(\out[1546]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [558]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[558]_i_2 
       (.I0(\f_permutation_l_/round_in [1226]),
        .I1(\f_permutation_l_/round_in [1290]),
        .I2(\out[1546]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[558]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[559]_i_1 
       (.I0(\out[559]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[869] ),
        .I2(\out[1553]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[480] ),
        .I4(\out[1547]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [559]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[559]_i_2 
       (.I0(\f_permutation_l_/round_in [1227]),
        .I1(\f_permutation_l_/round_in [1291]),
        .I2(\out[1547]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[559]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[55]_i_1 
       (.I0(\out[1569]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[245] ),
        .I2(\out[311]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1024]),
        .I4(\out[1493]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[560]_i_1 
       (.I0(\out[560]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[870] ),
        .I2(\out[1554]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[481] ),
        .I4(\out[1548]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [560]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[560]_i_2 
       (.I0(\f_permutation_l_/round_in [1228]),
        .I1(\f_permutation_l_/round_in [1292]),
        .I2(\out[1548]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[560]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[561]_i_1 
       (.I0(\out[561]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[871] ),
        .I2(\out[1555]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[482] ),
        .I4(\out[1549]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [561]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[561]_i_2 
       (.I0(\f_permutation_l_/round_in [1229]),
        .I1(\f_permutation_l_/round_in [1293]),
        .I2(\out[1549]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[561]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[562]_i_1 
       (.I0(\out[562]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[872] ),
        .I2(\out[1556]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[483] ),
        .I4(\out[1550]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [562]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[562]_i_2 
       (.I0(\f_permutation_l_/round_in [1230]),
        .I1(\f_permutation_l_/round_in [1294]),
        .I2(\out[1550]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[562]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[563]_i_1 
       (.I0(\out[563]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[873] ),
        .I2(\out[1557]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[484] ),
        .I4(\out[1551]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [563]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[563]_i_2 
       (.I0(\f_permutation_l_/round_in [1231]),
        .I1(\f_permutation_l_/round_in [1295]),
        .I2(\out[1551]_i_15_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[563]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[564]_i_1 
       (.I0(\out[564]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[874] ),
        .I2(\out[1558]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[485] ),
        .I4(\out[1552]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [564]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[564]_i_2 
       (.I0(\f_permutation_l_/round_in [1232]),
        .I1(\f_permutation_l_/round_in [1296]),
        .I2(\out[1552]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[564]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[565]_i_1 
       (.I0(\out[565]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[875] ),
        .I2(\out[1559]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[486] ),
        .I4(\out[1553]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [565]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[565]_i_2 
       (.I0(\f_permutation_l_/round_in [1233]),
        .I1(\f_permutation_l_/round_in [1297]),
        .I2(\out[1553]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[565]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[566]_i_1 
       (.I0(\out[566]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[876] ),
        .I2(\out[1560]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[487] ),
        .I4(\out[1554]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [566]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[566]_i_2 
       (.I0(\f_permutation_l_/round_in [1234]),
        .I1(\f_permutation_l_/round_in [1298]),
        .I2(\out[1554]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[566]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[567]_i_1 
       (.I0(\out[567]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[877] ),
        .I2(\out[1561]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[488] ),
        .I4(\out[1555]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [567]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[567]_i_2 
       (.I0(\f_permutation_l_/round_in [1235]),
        .I1(\f_permutation_l_/round_in [1299]),
        .I2(\out[1555]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[567]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[568]_i_1 
       (.I0(\out[568]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[878] ),
        .I2(\out[1562]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[489] ),
        .I4(\out[1556]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [568]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[568]_i_2 
       (.I0(\f_permutation_l_/round_in [1236]),
        .I1(\f_permutation_l_/round_in [1300]),
        .I2(\out[1556]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[568]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[569]_i_1 
       (.I0(\out[569]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[879] ),
        .I2(\out[1563]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[490] ),
        .I4(\out[1557]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [569]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[569]_i_2 
       (.I0(\f_permutation_l_/round_in [1237]),
        .I1(\f_permutation_l_/round_in [1301]),
        .I2(\out[1557]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[569]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[56]_i_1 
       (.I0(\out[1570]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[246] ),
        .I2(\out[312]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1025]),
        .I4(\out[1494]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[570]_i_1 
       (.I0(\out[570]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[880] ),
        .I2(\out[1564]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[491] ),
        .I4(\out[1558]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [570]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[570]_i_2 
       (.I0(\f_permutation_l_/round_in [1238]),
        .I1(\out[1536]_i_14_n_0 ),
        .I2(\f_permutation_l_/round_in [1493]),
        .I3(\f_permutation_l_/round_in [1302]),
        .I4(\out[1558]_i_14_n_0 ),
        .O(\out[570]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[571]_i_1 
       (.I0(\out[571]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[881] ),
        .I2(\out[1565]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[492] ),
        .I4(\out[1559]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [571]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[571]_i_2 
       (.I0(\f_permutation_l_/round_in [1239]),
        .I1(\f_permutation_l_/round_in [1494]),
        .I2(\out[1537]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1303]),
        .I4(\out[1559]_i_15_n_0 ),
        .O(\out[571]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[572]_i_1 
       (.I0(\out[572]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[882] ),
        .I2(\out[1566]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[493] ),
        .I4(\out[1560]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [572]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[572]_i_2 
       (.I0(\f_permutation_l_/round_in [1240]),
        .I1(\f_permutation_l_/round_in [1495]),
        .I2(\out[1538]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1304]),
        .I4(\out[1560]_i_15_n_0 ),
        .O(\out[572]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[573]_i_1 
       (.I0(\out[573]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[883] ),
        .I2(\out[1311]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[494] ),
        .I4(\out[1561]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [573]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[573]_i_2 
       (.I0(\f_permutation_l_/round_in [1241]),
        .I1(\f_permutation_l_/round_in [1496]),
        .I2(\out[1539]_i_14_n_0 ),
        .I3(\f_permutation_l_/round_in [1305]),
        .I4(\out[1561]_i_14_n_0 ),
        .O(\out[573]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[574]_i_1 
       (.I0(\out[574]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[884] ),
        .I2(\out[1568]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[495] ),
        .I4(\out[1562]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [574]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[574]_i_2 
       (.I0(\f_permutation_l_/round_in [1242]),
        .I1(\f_permutation_l_/round_in [1497]),
        .I2(\out[1540]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1306]),
        .I4(\out[1562]_i_15_n_0 ),
        .O(\out[574]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69AAAA69)) 
    \out[575]_i_1 
       (.I0(\out[575]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[885] ),
        .I2(\out[1569]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[496] ),
        .I4(\out[1563]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [575]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[575]_i_2 
       (.I0(\f_permutation_l_/round_in [1243]),
        .I1(\f_permutation_l_/round_in [1498]),
        .I2(\out[1541]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1307]),
        .I4(\out[1563]_i_14_n_0 ),
        .O(\out[575]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[576]_i_1 
       (.I0(\f_permutation_l_/round_in [1244]),
        .I1(\out[1247]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[886] ),
        .I3(\out[1570]_i_3_n_0 ),
        .I4(\out[576]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [576]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[576]_i_2 
       (.I0(padder_out_1[228]),
        .I1(out[164]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1244]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[576]_i_3 
       (.I0(\f_permutation_l_/round_in [1317]),
        .I1(\out[1552]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1572]),
        .I3(\f_permutation_l_/round_in [1381]),
        .I4(\out[1553]_i_10_n_0 ),
        .O(\out[576]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[577]_i_1 
       (.I0(\f_permutation_l_/round_in [1245]),
        .I1(\out[1248]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[887] ),
        .I3(\out[1571]_i_3_n_0 ),
        .I4(\out[577]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [577]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[577]_i_2 
       (.I0(padder_out_1[229]),
        .I1(out[165]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1245]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[577]_i_3 
       (.I0(\f_permutation_l_/round_in [1318]),
        .I1(\out[1553]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1573]),
        .I3(\f_permutation_l_/round_in [1382]),
        .I4(\out[1554]_i_10_n_0 ),
        .O(\out[577]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[578]_i_1 
       (.I0(\f_permutation_l_/round_in [1246]),
        .I1(\out[1249]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[888] ),
        .I3(\out[1572]_i_3_n_0 ),
        .I4(\out[578]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [578]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[578]_i_2 
       (.I0(padder_out_1[230]),
        .I1(out[166]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1246]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[578]_i_3 
       (.I0(\f_permutation_l_/round_in [1319]),
        .I1(\out[1554]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1574]),
        .I3(\f_permutation_l_/round_in [1383]),
        .I4(\out[1555]_i_10_n_0 ),
        .O(\out[578]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[579]_i_1 
       (.I0(\f_permutation_l_/round_in [1247]),
        .I1(\out[1250]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[889] ),
        .I3(\out[1573]_i_3_n_0 ),
        .I4(\out[579]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [579]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[579]_i_2 
       (.I0(padder_out_1[231]),
        .I1(out[167]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1247]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[579]_i_3 
       (.I0(\f_permutation_l_/round_in [1320]),
        .I1(\out[1555]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1575]),
        .I3(\f_permutation_l_/round_in [1384]),
        .I4(\out[1556]_i_11_n_0 ),
        .O(\out[579]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[57]_i_1 
       (.I0(\out[1571]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[247] ),
        .I2(\out[313]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1026]),
        .I4(\out[1495]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[580]_i_1 
       (.I0(\f_permutation_l_/round_in [1248]),
        .I1(\out[1251]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[890] ),
        .I3(\out[1574]_i_3_n_0 ),
        .I4(\out[580]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [580]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[580]_i_2 
       (.I0(padder_out_1[216]),
        .I1(out[152]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1248]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[580]_i_3 
       (.I0(\f_permutation_l_/round_in [1321]),
        .I1(\out[1556]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1576]),
        .I3(\f_permutation_l_/round_in [1385]),
        .I4(\out[1557]_i_10_n_0 ),
        .O(\out[580]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[581]_i_1 
       (.I0(\f_permutation_l_/round_in [1249]),
        .I1(\out[1252]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[891] ),
        .I3(\out[1575]_i_3_n_0 ),
        .I4(\out[581]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [581]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[581]_i_2 
       (.I0(padder_out_1[217]),
        .I1(out[153]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1249]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[581]_i_3 
       (.I0(\f_permutation_l_/round_in [1322]),
        .I1(\out[1557]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1577]),
        .I3(\f_permutation_l_/round_in [1386]),
        .I4(\out[1558]_i_10_n_0 ),
        .O(\out[581]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[582]_i_1 
       (.I0(\f_permutation_l_/round_in [1250]),
        .I1(\out[1253]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[892] ),
        .I3(\out[1576]_i_3_n_0 ),
        .I4(\out[582]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [582]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[582]_i_2 
       (.I0(padder_out_1[218]),
        .I1(out[154]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1250]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[582]_i_3 
       (.I0(\f_permutation_l_/round_in [1323]),
        .I1(\out[1558]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1578]),
        .I3(\f_permutation_l_/round_in [1387]),
        .I4(\out[1559]_i_10_n_0 ),
        .O(\out[582]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[583]_i_1 
       (.I0(\f_permutation_l_/round_in [1251]),
        .I1(\out[1254]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[893] ),
        .I3(\out[1577]_i_3_n_0 ),
        .I4(\out[583]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [583]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[583]_i_2 
       (.I0(padder_out_1[219]),
        .I1(out[155]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1251]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[583]_i_3 
       (.I0(\f_permutation_l_/round_in [1324]),
        .I1(\out[1559]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1579]),
        .I3(\f_permutation_l_/round_in [1388]),
        .I4(\out[1560]_i_10_n_0 ),
        .O(\out[583]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[584]_i_1 
       (.I0(\f_permutation_l_/round_in [1252]),
        .I1(\out[1255]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[894] ),
        .I3(\out[1578]_i_3_n_0 ),
        .I4(\out[584]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [584]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[584]_i_2 
       (.I0(padder_out_1[220]),
        .I1(out[156]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1252]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[584]_i_3 
       (.I0(\f_permutation_l_/round_in [1325]),
        .I1(\out[1560]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1580]),
        .I3(\f_permutation_l_/round_in [1389]),
        .I4(\out[1561]_i_10_n_0 ),
        .O(\out[584]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[585]_i_1 
       (.I0(\f_permutation_l_/round_in [1253]),
        .I1(\out[1256]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[895] ),
        .I3(\out[1579]_i_3_n_0 ),
        .I4(\out[585]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [585]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[585]_i_2 
       (.I0(padder_out_1[221]),
        .I1(out[157]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1253]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[585]_i_3 
       (.I0(\f_permutation_l_/round_in [1326]),
        .I1(\out[1561]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1581]),
        .I3(\f_permutation_l_/round_in [1390]),
        .I4(\out[1562]_i_10_n_0 ),
        .O(\out[585]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[586]_i_1 
       (.I0(\f_permutation_l_/round_in [1254]),
        .I1(\out[1257]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[832] ),
        .I3(\out[1580]_i_3_n_0 ),
        .I4(\out[586]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [586]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[586]_i_2 
       (.I0(padder_out_1[222]),
        .I1(out[158]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1254]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[586]_i_3 
       (.I0(\f_permutation_l_/round_in [1327]),
        .I1(\out[1562]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1582]),
        .I3(\f_permutation_l_/round_in [1391]),
        .I4(\out[1563]_i_10_n_0 ),
        .O(\out[586]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[587]_i_1 
       (.I0(\f_permutation_l_/round_in [1255]),
        .I1(\out[1258]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[833] ),
        .I3(\out[1581]_i_3_n_0 ),
        .I4(\out[587]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [587]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[587]_i_2 
       (.I0(padder_out_1[223]),
        .I1(out[159]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1255]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[587]_i_3 
       (.I0(\f_permutation_l_/round_in [1328]),
        .I1(\out[1563]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1583]),
        .I3(\f_permutation_l_/round_in [1392]),
        .I4(\out[1564]_i_10_n_0 ),
        .O(\out[587]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[588]_i_1 
       (.I0(\f_permutation_l_/round_in [1256]),
        .I1(\out[1259]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[834] ),
        .I3(\out[1582]_i_3_n_0 ),
        .I4(\out[588]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [588]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[588]_i_2 
       (.I0(padder_out_1[208]),
        .I1(out[144]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1256]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[588]_i_3 
       (.I0(\f_permutation_l_/round_in [1329]),
        .I1(\out[1564]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1584]),
        .I3(\f_permutation_l_/round_in [1393]),
        .I4(\out[1565]_i_10_n_0 ),
        .O(\out[588]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[589]_i_1 
       (.I0(\f_permutation_l_/round_in [1257]),
        .I1(\out[1260]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[835] ),
        .I3(\out[1583]_i_3_n_0 ),
        .I4(\out[589]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [589]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[589]_i_2 
       (.I0(padder_out_1[209]),
        .I1(out[145]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1257]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[589]_i_3 
       (.I0(\f_permutation_l_/round_in [1330]),
        .I1(\out[1565]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1585]),
        .I3(\f_permutation_l_/round_in [1394]),
        .I4(\out[1566]_i_10_n_0 ),
        .O(\out[589]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[58]_i_1 
       (.I0(\out[1572]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[248] ),
        .I2(\out[314]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1027]),
        .I4(\out[1496]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[590]_i_1 
       (.I0(\f_permutation_l_/round_in [1258]),
        .I1(\out[1261]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[836] ),
        .I3(\out[1584]_i_3_n_0 ),
        .I4(\out[590]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [590]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[590]_i_2 
       (.I0(padder_out_1[210]),
        .I1(out[146]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1258]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[590]_i_3 
       (.I0(\f_permutation_l_/round_in [1331]),
        .I1(\out[1566]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1586]),
        .I3(\f_permutation_l_/round_in [1395]),
        .I4(\out[1567]_i_11_n_0 ),
        .O(\out[590]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[591]_i_1 
       (.I0(\f_permutation_l_/round_in [1259]),
        .I1(\out[1262]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[837] ),
        .I3(\out[1585]_i_3_n_0 ),
        .I4(\out[591]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [591]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[591]_i_2 
       (.I0(padder_out_1[211]),
        .I1(out[147]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1259]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[591]_i_3 
       (.I0(\f_permutation_l_/round_in [1332]),
        .I1(\out[1567]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1587]),
        .I3(\f_permutation_l_/round_in [1396]),
        .I4(\out[1568]_i_10_n_0 ),
        .O(\out[591]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[592]_i_1 
       (.I0(\f_permutation_l_/round_in [1260]),
        .I1(\out[1263]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[838] ),
        .I3(\out[1586]_i_3_n_0 ),
        .I4(\out[592]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [592]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[592]_i_2 
       (.I0(padder_out_1[212]),
        .I1(out[148]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1260]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[592]_i_3 
       (.I0(\f_permutation_l_/round_in [1333]),
        .I1(\out[1568]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1588]),
        .I3(\f_permutation_l_/round_in [1397]),
        .I4(\out[1569]_i_10_n_0 ),
        .O(\out[592]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[593]_i_1 
       (.I0(\f_permutation_l_/round_in [1261]),
        .I1(\out[1264]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[839] ),
        .I3(\out[1587]_i_3_n_0 ),
        .I4(\out[593]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [593]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[593]_i_2 
       (.I0(padder_out_1[213]),
        .I1(out[149]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1261]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[593]_i_3 
       (.I0(\f_permutation_l_/round_in [1334]),
        .I1(\out[1569]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1589]),
        .I3(\f_permutation_l_/round_in [1398]),
        .I4(\out[1570]_i_10_n_0 ),
        .O(\out[593]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[594]_i_1 
       (.I0(\f_permutation_l_/round_in [1262]),
        .I1(\out[1265]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[840] ),
        .I3(\out[1588]_i_3_n_0 ),
        .I4(\out[594]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [594]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[594]_i_2 
       (.I0(padder_out_1[214]),
        .I1(out[150]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1262]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[594]_i_3 
       (.I0(\f_permutation_l_/round_in [1335]),
        .I1(\out[1570]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1590]),
        .I3(\f_permutation_l_/round_in [1399]),
        .I4(\out[1571]_i_10_n_0 ),
        .O(\out[594]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[595]_i_1 
       (.I0(\f_permutation_l_/round_in [1263]),
        .I1(\out[1266]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[841] ),
        .I3(\out[1589]_i_3_n_0 ),
        .I4(\out[595]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [595]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[595]_i_2 
       (.I0(padder_out_1[215]),
        .I1(out[151]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1263]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[595]_i_3 
       (.I0(\f_permutation_l_/round_in [1336]),
        .I1(\out[1571]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1591]),
        .I3(\f_permutation_l_/round_in [1400]),
        .I4(\out[1572]_i_10_n_0 ),
        .O(\out[595]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[596]_i_1 
       (.I0(\f_permutation_l_/round_in [1264]),
        .I1(\out[1267]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[842] ),
        .I3(\out[1590]_i_3_n_0 ),
        .I4(\out[596]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [596]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[596]_i_2 
       (.I0(padder_out_1[200]),
        .I1(out[136]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1264]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[596]_i_3 
       (.I0(\f_permutation_l_/round_in [1337]),
        .I1(\out[1572]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1592]),
        .I3(\f_permutation_l_/round_in [1401]),
        .I4(\out[1573]_i_10_n_0 ),
        .O(\out[596]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[597]_i_1 
       (.I0(\f_permutation_l_/round_in [1265]),
        .I1(\out[1268]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[843] ),
        .I3(\out[1591]_i_3_n_0 ),
        .I4(\out[597]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [597]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[597]_i_2 
       (.I0(padder_out_1[201]),
        .I1(out[137]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1265]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[597]_i_3 
       (.I0(\f_permutation_l_/round_in [1338]),
        .I1(\out[1573]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1593]),
        .I3(\f_permutation_l_/round_in [1402]),
        .I4(\out[1574]_i_10_n_0 ),
        .O(\out[597]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[598]_i_1 
       (.I0(\f_permutation_l_/round_in [1266]),
        .I1(\out[1269]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[844] ),
        .I3(\out[1592]_i_3_n_0 ),
        .I4(\out[598]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [598]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[598]_i_2 
       (.I0(padder_out_1[202]),
        .I1(out[138]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1266]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[598]_i_3 
       (.I0(\f_permutation_l_/round_in [1339]),
        .I1(\out[1574]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1594]),
        .I3(\f_permutation_l_/round_in [1403]),
        .I4(\out[1575]_i_10_n_0 ),
        .O(\out[598]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[599]_i_1 
       (.I0(\f_permutation_l_/round_in [1267]),
        .I1(\out[1270]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[845] ),
        .I3(\out[1593]_i_3_n_0 ),
        .I4(\out[599]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [599]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[599]_i_2 
       (.I0(padder_out_1[203]),
        .I1(out[139]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1267]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[599]_i_3 
       (.I0(\f_permutation_l_/round_in [1340]),
        .I1(\out[1575]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1595]),
        .I3(\f_permutation_l_/round_in [1404]),
        .I4(\out[1576]_i_10_n_0 ),
        .O(\out[599]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[59]_i_1 
       (.I0(\out[1573]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[249] ),
        .I2(\out[315]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1028]),
        .I4(\out[1497]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[5]_i_1 
       (.I0(\out[1583]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[195] ),
        .I2(\out[261]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1038]),
        .I4(\out[1507]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[600]_i_1 
       (.I0(\f_permutation_l_/round_in [1268]),
        .I1(\out[1271]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[846] ),
        .I3(\out[1594]_i_3_n_0 ),
        .I4(\out[600]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [600]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[600]_i_2 
       (.I0(padder_out_1[204]),
        .I1(out[140]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1268]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[600]_i_3 
       (.I0(\f_permutation_l_/round_in [1341]),
        .I1(\out[1576]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1596]),
        .I3(\f_permutation_l_/round_in [1405]),
        .I4(\out[1577]_i_10_n_0 ),
        .O(\out[600]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[601]_i_1 
       (.I0(\f_permutation_l_/round_in [1269]),
        .I1(\out[1272]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[847] ),
        .I3(\out[1595]_i_3_n_0 ),
        .I4(\out[601]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [601]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[601]_i_2 
       (.I0(padder_out_1[205]),
        .I1(out[141]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1269]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[601]_i_3 
       (.I0(\f_permutation_l_/round_in [1342]),
        .I1(\f_permutation_l_/round_in [1597]),
        .I2(\out[1577]_i_6_n_0 ),
        .I3(\out[1578]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1406]),
        .O(\out[601]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[602]_i_1 
       (.I0(\f_permutation_l_/round_in [1270]),
        .I1(\out[1273]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[848] ),
        .I3(\out[1596]_i_3_n_0 ),
        .I4(\out[602]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [602]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[602]_i_2 
       (.I0(padder_out_1[206]),
        .I1(out[142]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1270]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[602]_i_3 
       (.I0(\f_permutation_l_/round_in [1343]),
        .I1(\f_permutation_l_/round_in [1598]),
        .I2(\out[1578]_i_6_n_0 ),
        .I3(\out[1579]_i_10_n_0 ),
        .I4(\f_permutation_l_/round_in [1407]),
        .O(\out[602]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[603]_i_1 
       (.I0(\f_permutation_l_/round_in [1271]),
        .I1(\out[1274]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[849] ),
        .I3(\out[1597]_i_3_n_0 ),
        .I4(\out[603]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [603]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[603]_i_2 
       (.I0(padder_out_1[207]),
        .I1(out[143]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1271]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[603]_i_3 
       (.I0(\f_permutation_l_/round_in [1280]),
        .I1(\f_permutation_l_/round_in [1599]),
        .I2(\out[1579]_i_7_n_0 ),
        .I3(\out[1580]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1344]),
        .O(\out[603]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[604]_i_1 
       (.I0(\f_permutation_l_/round_in [1272]),
        .I1(\out[1275]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[850] ),
        .I3(\out[1598]_i_3_n_0 ),
        .I4(\out[604]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [604]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[604]_i_2 
       (.I0(padder_out_1[192]),
        .I1(out[128]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1272]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[604]_i_3 
       (.I0(\f_permutation_l_/round_in [1281]),
        .I1(\f_permutation_l_/round_in [1536]),
        .I2(\out[1580]_i_6_n_0 ),
        .I3(\out[1581]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1345]),
        .O(\out[604]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[605]_i_1 
       (.I0(\f_permutation_l_/round_in [1273]),
        .I1(\out[1276]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[851] ),
        .I3(\out[1343]_i_3_n_0 ),
        .I4(\out[605]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [605]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[605]_i_2 
       (.I0(padder_out_1[193]),
        .I1(out[129]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1273]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[605]_i_3 
       (.I0(\f_permutation_l_/round_in [1282]),
        .I1(\f_permutation_l_/round_in [1537]),
        .I2(\out[1581]_i_6_n_0 ),
        .I3(\out[1582]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1346]),
        .O(\out[605]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[606]_i_1 
       (.I0(\f_permutation_l_/round_in [1274]),
        .I1(\out[1277]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[852] ),
        .I3(\out[1280]_i_3_n_0 ),
        .I4(\out[606]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [606]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[606]_i_2 
       (.I0(padder_out_1[194]),
        .I1(out[130]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1274]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[606]_i_3 
       (.I0(\f_permutation_l_/round_in [1283]),
        .I1(\f_permutation_l_/round_in [1538]),
        .I2(\out[1582]_i_6_n_0 ),
        .I3(\out[1583]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1347]),
        .O(\out[606]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[607]_i_1 
       (.I0(\f_permutation_l_/round_in [1275]),
        .I1(\out[1278]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[853] ),
        .I3(\out[1281]_i_3_n_0 ),
        .I4(\out[607]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [607]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[607]_i_2 
       (.I0(padder_out_1[195]),
        .I1(out[131]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1275]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[607]_i_3 
       (.I0(\f_permutation_l_/round_in [1284]),
        .I1(\f_permutation_l_/round_in [1539]),
        .I2(\out[1583]_i_6_n_0 ),
        .I3(\out[1584]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1348]),
        .O(\out[607]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[608]_i_1 
       (.I0(\f_permutation_l_/round_in [1276]),
        .I1(\out[1279]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[854] ),
        .I3(\out[1538]_i_3_n_0 ),
        .I4(\out[608]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [608]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[608]_i_2 
       (.I0(padder_out_1[196]),
        .I1(out[132]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1276]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[608]_i_3 
       (.I0(\f_permutation_l_/round_in [1285]),
        .I1(\f_permutation_l_/round_in [1540]),
        .I2(\out[1584]_i_6_n_0 ),
        .I3(\out[1585]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1349]),
        .O(\out[608]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[609]_i_1 
       (.I0(\f_permutation_l_/round_in [1277]),
        .I1(\out[1216]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[855] ),
        .I3(\out[1539]_i_3_n_0 ),
        .I4(\out[609]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [609]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[609]_i_2 
       (.I0(padder_out_1[197]),
        .I1(out[133]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1277]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[609]_i_3 
       (.I0(\f_permutation_l_/round_in [1286]),
        .I1(\f_permutation_l_/round_in [1541]),
        .I2(\out[1585]_i_6_n_0 ),
        .I3(\out[1586]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1350]),
        .O(\out[609]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[60]_i_1 
       (.I0(\out[1574]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[250] ),
        .I2(\out[316]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1029]),
        .I4(\out[1498]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[610]_i_1 
       (.I0(\f_permutation_l_/round_in [1278]),
        .I1(\out[1217]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[856] ),
        .I3(\out[1540]_i_3_n_0 ),
        .I4(\out[610]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [610]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[610]_i_2 
       (.I0(padder_out_1[198]),
        .I1(out[134]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1278]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[610]_i_3 
       (.I0(\f_permutation_l_/round_in [1287]),
        .I1(\f_permutation_l_/round_in [1542]),
        .I2(\out[1586]_i_6_n_0 ),
        .I3(\out[1587]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1351]),
        .O(\out[610]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[611]_i_1 
       (.I0(\f_permutation_l_/round_in [1279]),
        .I1(\out[1218]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[857] ),
        .I3(\out[1541]_i_3_n_0 ),
        .I4(\out[611]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [611]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[611]_i_2 
       (.I0(padder_out_1[199]),
        .I1(out[135]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1279]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[611]_i_3 
       (.I0(\f_permutation_l_/round_in [1288]),
        .I1(\f_permutation_l_/round_in [1543]),
        .I2(\out[1587]_i_6_n_0 ),
        .I3(\out[1588]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1352]),
        .O(\out[611]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[612]_i_1 
       (.I0(\f_permutation_l_/round_in [1216]),
        .I1(\out[1219]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[858] ),
        .I3(\out[1542]_i_3_n_0 ),
        .I4(\out[612]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [612]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[612]_i_2 
       (.I0(padder_out_1[248]),
        .I1(out[184]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1216]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[612]_i_3 
       (.I0(\f_permutation_l_/round_in [1289]),
        .I1(\f_permutation_l_/round_in [1544]),
        .I2(\out[1588]_i_6_n_0 ),
        .I3(\out[1589]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1353]),
        .O(\out[612]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[613]_i_1 
       (.I0(\f_permutation_l_/round_in [1217]),
        .I1(\out[1220]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[859] ),
        .I3(\out[1287]_i_3_n_0 ),
        .I4(\out[613]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [613]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[613]_i_2 
       (.I0(padder_out_1[249]),
        .I1(out[185]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1217]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[613]_i_3 
       (.I0(\f_permutation_l_/round_in [1290]),
        .I1(\f_permutation_l_/round_in [1545]),
        .I2(\out[1589]_i_6_n_0 ),
        .I3(\out[1590]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1354]),
        .O(\out[613]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[614]_i_1 
       (.I0(\f_permutation_l_/round_in [1218]),
        .I1(\out[1221]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[860] ),
        .I3(\out[1544]_i_3_n_0 ),
        .I4(\out[614]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [614]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[614]_i_2 
       (.I0(padder_out_1[250]),
        .I1(out[186]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1218]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[614]_i_3 
       (.I0(\f_permutation_l_/round_in [1291]),
        .I1(\f_permutation_l_/round_in [1546]),
        .I2(\out[1590]_i_6_n_0 ),
        .I3(\out[1591]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1355]),
        .O(\out[614]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[615]_i_1 
       (.I0(\f_permutation_l_/round_in [1219]),
        .I1(\out[1539]_i_6_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[861] ),
        .I3(\out[1545]_i_3_n_0 ),
        .I4(\out[615]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [615]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[615]_i_2 
       (.I0(padder_out_1[251]),
        .I1(out[187]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1219]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[615]_i_3 
       (.I0(\f_permutation_l_/round_in [1292]),
        .I1(\f_permutation_l_/round_in [1547]),
        .I2(\out[1591]_i_6_n_0 ),
        .I3(\out[1592]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1356]),
        .O(\out[615]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[616]_i_1 
       (.I0(\f_permutation_l_/round_in [1220]),
        .I1(\out[1223]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[862] ),
        .I3(\out[1546]_i_3_n_0 ),
        .I4(\out[616]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [616]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[616]_i_2 
       (.I0(padder_out_1[252]),
        .I1(out[188]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1220]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[616]_i_3 
       (.I0(\f_permutation_l_/round_in [1293]),
        .I1(\f_permutation_l_/round_in [1548]),
        .I2(\out[1592]_i_6_n_0 ),
        .I3(\out[1593]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1357]),
        .O(\out[616]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[617]_i_1 
       (.I0(\f_permutation_l_/round_in [1221]),
        .I1(\out[1224]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[863] ),
        .I3(\out[1547]_i_3_n_0 ),
        .I4(\out[617]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [617]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[617]_i_2 
       (.I0(padder_out_1[253]),
        .I1(out[189]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1221]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[617]_i_3 
       (.I0(\f_permutation_l_/round_in [1294]),
        .I1(\f_permutation_l_/round_in [1549]),
        .I2(\out[1593]_i_6_n_0 ),
        .I3(\out[1594]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1358]),
        .O(\out[617]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[618]_i_1 
       (.I0(\f_permutation_l_/round_in [1222]),
        .I1(\out[1225]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[864] ),
        .I3(\out[1548]_i_3_n_0 ),
        .I4(\out[618]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [618]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[618]_i_2 
       (.I0(padder_out_1[254]),
        .I1(out[190]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1222]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[618]_i_3 
       (.I0(\f_permutation_l_/round_in [1295]),
        .I1(\f_permutation_l_/round_in [1550]),
        .I2(\out[1594]_i_6_n_0 ),
        .I3(\out[1595]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1359]),
        .O(\out[618]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[619]_i_1 
       (.I0(\f_permutation_l_/round_in [1223]),
        .I1(\out[1226]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[865] ),
        .I3(\out[1549]_i_3_n_0 ),
        .I4(\out[619]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [619]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[619]_i_2 
       (.I0(padder_out_1[255]),
        .I1(out[191]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1223]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[619]_i_3 
       (.I0(\f_permutation_l_/round_in [1296]),
        .I1(\f_permutation_l_/round_in [1551]),
        .I2(\out[1595]_i_6_n_0 ),
        .I3(\out[1596]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1360]),
        .O(\out[619]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[61]_i_1 
       (.I0(\out[1575]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[251] ),
        .I2(\out[317]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1030]),
        .I4(\out[1499]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[620]_i_1 
       (.I0(\f_permutation_l_/round_in [1224]),
        .I1(\out[1227]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[866] ),
        .I3(\out[1550]_i_3_n_0 ),
        .I4(\out[620]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [620]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[620]_i_2 
       (.I0(padder_out_1[240]),
        .I1(out[176]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1224]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[620]_i_3 
       (.I0(\f_permutation_l_/round_in [1297]),
        .I1(\f_permutation_l_/round_in [1552]),
        .I2(\out[1596]_i_6_n_0 ),
        .I3(\out[1597]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1361]),
        .O(\out[620]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[621]_i_1 
       (.I0(\f_permutation_l_/round_in [1225]),
        .I1(\out[1228]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[867] ),
        .I3(\out[1295]_i_3_n_0 ),
        .I4(\out[621]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [621]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[621]_i_2 
       (.I0(padder_out_1[241]),
        .I1(out[177]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1225]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[621]_i_3 
       (.I0(\f_permutation_l_/round_in [1298]),
        .I1(\f_permutation_l_/round_in [1553]),
        .I2(\out[1597]_i_6_n_0 ),
        .I3(\out[1598]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1362]),
        .O(\out[621]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[622]_i_1 
       (.I0(\f_permutation_l_/round_in [1226]),
        .I1(\out[1229]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[868] ),
        .I3(\out[1552]_i_3_n_0 ),
        .I4(\out[622]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [622]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[622]_i_2 
       (.I0(padder_out_1[242]),
        .I1(out[178]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1226]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[622]_i_3 
       (.I0(\f_permutation_l_/round_in [1299]),
        .I1(\f_permutation_l_/round_in [1554]),
        .I2(\out[1598]_i_6_n_0 ),
        .I3(\out[1599]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1363]),
        .O(\out[622]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[623]_i_1 
       (.I0(\f_permutation_l_/round_in [1227]),
        .I1(\out[1230]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[869] ),
        .I3(\out[1553]_i_3_n_0 ),
        .I4(\out[623]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [623]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[623]_i_2 
       (.I0(padder_out_1[243]),
        .I1(out[179]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1227]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[623]_i_3 
       (.I0(\f_permutation_l_/round_in [1300]),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1555]),
        .I4(\out[1599]_i_8_n_0 ),
        .O(\out[623]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[624]_i_1 
       (.I0(\f_permutation_l_/round_in [1228]),
        .I1(\out[1231]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[870] ),
        .I3(\out[1554]_i_3_n_0 ),
        .I4(\out[624]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [624]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[624]_i_2 
       (.I0(padder_out_1[244]),
        .I1(out[180]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1228]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[624]_i_3 
       (.I0(\f_permutation_l_/round_in [1301]),
        .I1(\out[1536]_i_10_n_0 ),
        .I2(\f_permutation_l_/round_in [1556]),
        .I3(\f_permutation_l_/round_in [1365]),
        .I4(\out[1537]_i_11_n_0 ),
        .O(\out[624]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[625]_i_1 
       (.I0(\f_permutation_l_/round_in [1229]),
        .I1(\out[1232]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[871] ),
        .I3(\out[1555]_i_3_n_0 ),
        .I4(\out[625]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [625]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[625]_i_2 
       (.I0(padder_out_1[245]),
        .I1(out[181]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1229]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[625]_i_3 
       (.I0(\f_permutation_l_/round_in [1302]),
        .I1(\out[1537]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1557]),
        .I3(\f_permutation_l_/round_in [1366]),
        .I4(\out[1538]_i_10_n_0 ),
        .O(\out[625]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[626]_i_1 
       (.I0(\f_permutation_l_/round_in [1230]),
        .I1(\out[1233]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[872] ),
        .I3(\out[1556]_i_3_n_0 ),
        .I4(\out[626]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [626]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[626]_i_2 
       (.I0(padder_out_1[246]),
        .I1(out[182]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1230]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[626]_i_3 
       (.I0(\f_permutation_l_/round_in [1303]),
        .I1(\f_permutation_l_/round_in [1558]),
        .I2(\out[1538]_i_6_n_0 ),
        .I3(\out[1539]_i_12_n_0 ),
        .I4(\f_permutation_l_/round_in [1367]),
        .O(\out[626]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[627]_i_1 
       (.I0(\f_permutation_l_/round_in [1231]),
        .I1(\out[1234]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[873] ),
        .I3(\out[1557]_i_3_n_0 ),
        .I4(\out[627]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [627]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[627]_i_2 
       (.I0(padder_out_1[247]),
        .I1(out[183]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1231]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[627]_i_3 
       (.I0(\f_permutation_l_/round_in [1304]),
        .I1(\out[1539]_i_8_n_0 ),
        .I2(\f_permutation_l_/round_in [1559]),
        .I3(\f_permutation_l_/round_in [1368]),
        .I4(\out[1540]_i_10_n_0 ),
        .O(\out[627]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[628]_i_1 
       (.I0(\f_permutation_l_/round_in [1232]),
        .I1(\out[1235]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[874] ),
        .I3(\out[1558]_i_3_n_0 ),
        .I4(\out[628]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [628]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[628]_i_2 
       (.I0(padder_out_1[232]),
        .I1(out[168]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1232]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[628]_i_3 
       (.I0(\f_permutation_l_/round_in [1305]),
        .I1(\out[1540]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1560]),
        .I3(\f_permutation_l_/round_in [1369]),
        .I4(\out[1541]_i_10_n_0 ),
        .O(\out[628]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[629]_i_1 
       (.I0(\f_permutation_l_/round_in [1233]),
        .I1(\out[1236]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[875] ),
        .I3(\out[1559]_i_3_n_0 ),
        .I4(\out[629]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [629]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[629]_i_2 
       (.I0(padder_out_1[233]),
        .I1(out[169]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1233]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[629]_i_3 
       (.I0(\f_permutation_l_/round_in [1306]),
        .I1(\out[1541]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1561]),
        .I3(\f_permutation_l_/round_in [1370]),
        .I4(\out[1542]_i_12_n_0 ),
        .O(\out[629]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[62]_i_1 
       (.I0(\out[1576]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[252] ),
        .I2(\out[318]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1031]),
        .I4(\out[1500]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[630]_i_1 
       (.I0(\f_permutation_l_/round_in [1234]),
        .I1(\out[1237]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[876] ),
        .I3(\out[1560]_i_3_n_0 ),
        .I4(\out[630]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [630]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[630]_i_2 
       (.I0(padder_out_1[234]),
        .I1(out[170]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1234]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[630]_i_3 
       (.I0(\f_permutation_l_/round_in [1307]),
        .I1(\out[1542]_i_7_n_0 ),
        .I2(\f_permutation_l_/round_in [1562]),
        .I3(\f_permutation_l_/round_in [1371]),
        .I4(\out[1543]_i_13_n_0 ),
        .O(\out[630]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[631]_i_1 
       (.I0(\f_permutation_l_/round_in [1235]),
        .I1(\out[1238]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[877] ),
        .I3(\out[1561]_i_3_n_0 ),
        .I4(\out[631]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [631]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[631]_i_2 
       (.I0(padder_out_1[235]),
        .I1(out[171]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1235]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[631]_i_3 
       (.I0(\f_permutation_l_/round_in [1308]),
        .I1(\out[1543]_i_10_n_0 ),
        .I2(\f_permutation_l_/round_in [1563]),
        .I3(\f_permutation_l_/round_in [1372]),
        .I4(\out[1544]_i_10_n_0 ),
        .O(\out[631]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[632]_i_1 
       (.I0(\f_permutation_l_/round_in [1236]),
        .I1(\out[1239]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[878] ),
        .I3(\out[1562]_i_3_n_0 ),
        .I4(\out[632]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [632]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[632]_i_2 
       (.I0(padder_out_1[236]),
        .I1(out[172]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1236]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[632]_i_3 
       (.I0(\f_permutation_l_/round_in [1309]),
        .I1(\out[1544]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1564]),
        .I3(\f_permutation_l_/round_in [1373]),
        .I4(\out[1545]_i_10_n_0 ),
        .O(\out[632]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[633]_i_1 
       (.I0(\f_permutation_l_/round_in [1237]),
        .I1(\out[1240]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[879] ),
        .I3(\out[1563]_i_3_n_0 ),
        .I4(\out[633]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [633]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[633]_i_2 
       (.I0(padder_out_1[237]),
        .I1(out[173]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1237]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[633]_i_3 
       (.I0(\f_permutation_l_/round_in [1310]),
        .I1(\out[1545]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1565]),
        .I3(\f_permutation_l_/round_in [1374]),
        .I4(\out[1546]_i_10_n_0 ),
        .O(\out[633]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF66F0990)) 
    \out[634]_i_1 
       (.I0(\f_permutation_l_/round_in [1238]),
        .I1(\out[1241]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[880] ),
        .I3(\out[1564]_i_3_n_0 ),
        .I4(\out[634]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [634]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[634]_i_2 
       (.I0(padder_out_1[238]),
        .I1(out[174]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1238]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[634]_i_3 
       (.I0(\f_permutation_l_/round_in [1311]),
        .I1(\out[1546]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1566]),
        .I3(\f_permutation_l_/round_in [1375]),
        .I4(\out[1547]_i_10_n_0 ),
        .O(\out[634]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[635]_i_1 
       (.I0(\f_permutation_l_/round_in [1239]),
        .I1(\out[1242]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[881] ),
        .I3(\out[1565]_i_3_n_0 ),
        .I4(\out[635]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [635]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[635]_i_2 
       (.I0(padder_out_1[239]),
        .I1(out[175]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1239]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[635]_i_3 
       (.I0(\f_permutation_l_/round_in [1312]),
        .I1(\out[1547]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1567]),
        .I3(\f_permutation_l_/round_in [1376]),
        .I4(\out[1548]_i_10_n_0 ),
        .O(\out[635]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[636]_i_1 
       (.I0(\f_permutation_l_/round_in [1240]),
        .I1(\out[1243]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[882] ),
        .I3(\out[1566]_i_3_n_0 ),
        .I4(\out[636]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [636]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[636]_i_2 
       (.I0(padder_out_1[224]),
        .I1(out[160]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1240]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[636]_i_3 
       (.I0(\f_permutation_l_/round_in [1313]),
        .I1(\out[1548]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1568]),
        .I3(\f_permutation_l_/round_in [1377]),
        .I4(\out[1549]_i_10_n_0 ),
        .O(\out[636]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[637]_i_1 
       (.I0(\f_permutation_l_/round_in [1241]),
        .I1(\out[1244]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[883] ),
        .I3(\out[1311]_i_3_n_0 ),
        .I4(\out[637]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [637]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[637]_i_2 
       (.I0(padder_out_1[225]),
        .I1(out[161]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1241]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[637]_i_3 
       (.I0(\f_permutation_l_/round_in [1314]),
        .I1(\out[1549]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1569]),
        .I3(\f_permutation_l_/round_in [1378]),
        .I4(\out[1550]_i_10_n_0 ),
        .O(\out[637]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[638]_i_1 
       (.I0(\f_permutation_l_/round_in [1242]),
        .I1(\out[1245]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[884] ),
        .I3(\out[1568]_i_3_n_0 ),
        .I4(\out[638]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [638]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[638]_i_2 
       (.I0(padder_out_1[226]),
        .I1(out[162]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1242]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[638]_i_3 
       (.I0(\f_permutation_l_/round_in [1315]),
        .I1(\out[1550]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1570]),
        .I3(\f_permutation_l_/round_in [1379]),
        .I4(\out[1551]_i_11_n_0 ),
        .O(\out[638]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[639]_i_1 
       (.I0(\f_permutation_l_/round_in [1243]),
        .I1(\out[1246]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[885] ),
        .I3(\out[1569]_i_3_n_0 ),
        .I4(\out[639]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [639]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[639]_i_2 
       (.I0(padder_out_1[227]),
        .I1(out[163]),
        .I2(\out[1579]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1243]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[639]_i_3 
       (.I0(\f_permutation_l_/round_in [1316]),
        .I1(\out[1551]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1571]),
        .I3(\f_permutation_l_/round_in [1380]),
        .I4(\out[1552]_i_10_n_0 ),
        .O(\out[639]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[63]_i_1 
       (.I0(\out[1577]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[253] ),
        .I2(\out[319]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1032]),
        .I4(\out[1501]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[640]_i_1 
       (.I0(\out[1265]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[302] ),
        .I2(\out[896]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1146]),
        .I4(\out[1573]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [640]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[641]_i_1 
       (.I0(\out[1266]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[303] ),
        .I2(\out[897]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1147]),
        .I4(\out[1574]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [641]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[642]_i_1 
       (.I0(\out[1267]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[304] ),
        .I2(\out[898]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1148]),
        .I4(\out[1575]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [642]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[643]_i_1 
       (.I0(\out[1268]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[305] ),
        .I2(\out[899]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1149]),
        .I4(\out[1576]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [643]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[644]_i_1 
       (.I0(\out[1269]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[306] ),
        .I2(\out[900]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1150]),
        .I4(\out[1577]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [644]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[645]_i_1 
       (.I0(\out[1270]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[307] ),
        .I2(\out[901]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1151]),
        .I4(\out[1578]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [645]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[646]_i_1 
       (.I0(\out[1271]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[308] ),
        .I2(\out[902]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1088]),
        .I4(\out[1579]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [646]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[647]_i_1 
       (.I0(\out[1272]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[309] ),
        .I2(\out[903]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1089]),
        .I4(\out[1580]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [647]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[648]_i_1 
       (.I0(\out[1273]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[310] ),
        .I2(\out[904]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1090]),
        .I4(\out[1581]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [648]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[649]_i_1 
       (.I0(\out[1274]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[311] ),
        .I2(\out[905]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1091]),
        .I4(\out[1582]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [649]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[64]_i_1 
       (.I0(\out[1242]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[599] ),
        .I2(\f_permutation_l_/out_reg_n_0_[254] ),
        .I3(\out[1578]_i_3_n_0 ),
        .I4(\out[256]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [64]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[650]_i_1 
       (.I0(\out[1275]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[312] ),
        .I2(\out[906]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1092]),
        .I4(\out[1583]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [650]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[651]_i_1 
       (.I0(\out[1276]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[313] ),
        .I2(\out[907]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1093]),
        .I4(\out[1584]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [651]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[652]_i_1 
       (.I0(\out[1277]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[314] ),
        .I2(\out[908]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1094]),
        .I4(\out[1585]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [652]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[653]_i_1 
       (.I0(\out[1278]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[315] ),
        .I2(\out[909]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1095]),
        .I4(\out[1586]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [653]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[654]_i_1 
       (.I0(\out[1279]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[316] ),
        .I2(\out[910]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1096]),
        .I4(\out[1587]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [654]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[655]_i_1 
       (.I0(\out[1216]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[317] ),
        .I2(\out[911]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1097]),
        .I4(\out[1588]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [655]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[656]_i_1 
       (.I0(\out[1217]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[318] ),
        .I2(\out[912]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1098]),
        .I4(\out[1589]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [656]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[657]_i_1 
       (.I0(\out[1218]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[319] ),
        .I2(\out[913]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1099]),
        .I4(\out[1590]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [657]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[658]_i_1 
       (.I0(\out[1219]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[256] ),
        .I2(\out[914]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1100]),
        .I4(\out[1591]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [658]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[659]_i_1 
       (.I0(\out[1220]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[257] ),
        .I2(\out[915]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1101]),
        .I4(\out[1592]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [659]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[65]_i_1 
       (.I0(\out[1243]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[600] ),
        .I2(\f_permutation_l_/out_reg_n_0_[255] ),
        .I3(\out[1579]_i_3_n_0 ),
        .I4(\out[257]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [65]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[660]_i_1 
       (.I0(\out[1221]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[258] ),
        .I2(\out[916]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1102]),
        .I4(\out[1593]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [660]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[661]_i_1 
       (.I0(\out[1539]_i_6_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[259] ),
        .I2(\out[917]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1103]),
        .I4(\out[1594]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [661]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[662]_i_1 
       (.I0(\out[1223]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[260] ),
        .I2(\out[918]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1104]),
        .I4(\out[1595]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [662]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[663]_i_1 
       (.I0(\out[1224]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[261] ),
        .I2(\out[919]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1105]),
        .I4(\out[1596]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [663]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[664]_i_1 
       (.I0(\out[1225]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[262] ),
        .I2(\out[920]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1106]),
        .I4(\out[1597]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [664]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[665]_i_1 
       (.I0(\out[1226]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[263] ),
        .I2(\out[921]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1107]),
        .I4(\out[1598]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [665]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[666]_i_1 
       (.I0(\out[1227]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[264] ),
        .I2(\out[922]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1108]),
        .I4(\out[1599]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [666]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[667]_i_1 
       (.I0(\out[1228]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[265] ),
        .I2(\out[923]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1109]),
        .I4(\out[1472]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [667]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[668]_i_1 
       (.I0(\out[1229]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[266] ),
        .I2(\out[924]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1110]),
        .I4(\out[1537]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [668]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[669]_i_1 
       (.I0(\out[1230]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[267] ),
        .I2(\out[925]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1111]),
        .I4(\out[1538]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [669]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[66]_i_1 
       (.I0(\out[1244]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[601] ),
        .I2(\f_permutation_l_/out_reg_n_0_[192] ),
        .I3(\out[1580]_i_3_n_0 ),
        .I4(\out[258]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [66]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[670]_i_1 
       (.I0(\out[1231]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[268] ),
        .I2(\f_permutation_l_/round_in [1501]),
        .I3(\out[1545]_i_3_n_0 ),
        .I4(\out[926]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [670]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[671]_i_1 
       (.I0(\out[1232]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[269] ),
        .I2(\out[927]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1113]),
        .I4(\out[1540]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [671]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[672]_i_1 
       (.I0(\out[1233]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[270] ),
        .I2(\out[928]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1114]),
        .I4(\out[1541]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [672]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[673]_i_1 
       (.I0(\out[1234]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[271] ),
        .I2(\out[929]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1115]),
        .I4(\out[1542]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [673]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[674]_i_1 
       (.I0(\out[1235]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[272] ),
        .I2(\out[930]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1116]),
        .I4(\out[1543]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [674]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[675]_i_1 
       (.I0(\out[1236]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[273] ),
        .I2(\out[931]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1117]),
        .I4(\out[1544]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [675]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[676]_i_1 
       (.I0(\out[1237]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[274] ),
        .I2(\out[932]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1118]),
        .I4(\out[1545]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [676]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[677]_i_1 
       (.I0(\out[1238]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[275] ),
        .I2(\out[933]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1119]),
        .I4(\out[1546]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [677]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[678]_i_1 
       (.I0(\out[1239]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[276] ),
        .I2(\out[934]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1120]),
        .I4(\out[1547]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [678]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[679]_i_1 
       (.I0(\out[1240]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[277] ),
        .I2(\out[935]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1121]),
        .I4(\out[1548]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [679]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[67]_i_1 
       (.I0(\out[1245]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[602] ),
        .I2(\f_permutation_l_/out_reg_n_0_[193] ),
        .I3(\out[1581]_i_3_n_0 ),
        .I4(\out[259]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [67]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[680]_i_1 
       (.I0(\out[1241]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[278] ),
        .I2(\out[936]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1122]),
        .I4(\out[1549]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [680]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[681]_i_1 
       (.I0(\out[1242]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[279] ),
        .I2(\out[937]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1123]),
        .I4(\out[1550]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [681]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[682]_i_1 
       (.I0(\out[1243]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[280] ),
        .I2(\out[938]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1124]),
        .I4(\out[1551]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [682]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[683]_i_1 
       (.I0(\out[1244]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[281] ),
        .I2(\out[939]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1125]),
        .I4(\out[1552]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [683]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[684]_i_1 
       (.I0(\out[1245]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[282] ),
        .I2(\out[940]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1126]),
        .I4(\out[1553]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [684]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[685]_i_1 
       (.I0(\out[1246]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[283] ),
        .I2(\out[941]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1127]),
        .I4(\out[1554]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [685]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[686]_i_1 
       (.I0(\out[1247]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[284] ),
        .I2(\out[942]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1128]),
        .I4(\out[1555]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [686]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[687]_i_1 
       (.I0(\out[1248]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[285] ),
        .I2(\out[943]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1129]),
        .I4(\out[1556]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [687]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[688]_i_1 
       (.I0(\out[1249]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[286] ),
        .I2(\out[944]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1130]),
        .I4(\out[1557]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [688]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[689]_i_1 
       (.I0(\out[1250]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[287] ),
        .I2(\out[945]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1131]),
        .I4(\out[1558]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [689]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[68]_i_1 
       (.I0(\out[1246]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[603] ),
        .I2(\f_permutation_l_/out_reg_n_0_[194] ),
        .I3(\out[1582]_i_3_n_0 ),
        .I4(\out[260]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [68]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[690]_i_1 
       (.I0(\out[1251]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[288] ),
        .I2(\out[946]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1132]),
        .I4(\out[1559]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [690]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[691]_i_1 
       (.I0(\out[1252]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[289] ),
        .I2(\out[947]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1133]),
        .I4(\out[1560]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [691]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[692]_i_1 
       (.I0(\out[1253]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[290] ),
        .I2(\out[948]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1134]),
        .I4(\out[1561]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [692]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[693]_i_1 
       (.I0(\out[1254]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[291] ),
        .I2(\out[949]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1135]),
        .I4(\out[1562]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [693]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[694]_i_1 
       (.I0(\out[1255]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[292] ),
        .I2(\out[950]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1136]),
        .I4(\out[1563]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [694]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[695]_i_1 
       (.I0(\out[1256]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[293] ),
        .I2(\out[951]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1137]),
        .I4(\out[1564]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [695]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[696]_i_1 
       (.I0(\out[1257]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[294] ),
        .I2(\out[952]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1138]),
        .I4(\out[1565]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [696]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[697]_i_1 
       (.I0(\out[1258]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[295] ),
        .I2(\out[953]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1139]),
        .I4(\out[1566]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [697]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[698]_i_1 
       (.I0(\out[1259]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[296] ),
        .I2(\out[954]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1140]),
        .I4(\out[1567]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [698]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[699]_i_1 
       (.I0(\out[1260]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[297] ),
        .I2(\out[955]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1141]),
        .I4(\out[1568]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [699]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[69]_i_1 
       (.I0(\out[1247]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[604] ),
        .I2(\f_permutation_l_/out_reg_n_0_[195] ),
        .I3(\out[1583]_i_3_n_0 ),
        .I4(\out[261]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [69]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[6]_i_1 
       (.I0(\out[1584]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[196] ),
        .I2(\out[262]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1039]),
        .I4(\out[1508]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[700]_i_1 
       (.I0(\out[1261]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[298] ),
        .I2(\out[956]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1142]),
        .I4(\out[1569]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [700]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[701]_i_1 
       (.I0(\out[1262]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[299] ),
        .I2(\out[957]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1143]),
        .I4(\out[1570]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [701]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[702]_i_1 
       (.I0(\out[1263]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[300] ),
        .I2(\out[958]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1144]),
        .I4(\out[1571]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [702]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[703]_i_1 
       (.I0(\out[1264]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[301] ),
        .I2(\out[959]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1145]),
        .I4(\out[1572]_i_4_n_0 ),
        .O(\f_permutation_l_/round_out [703]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[704]_i_1 
       (.I0(\out[1414]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[376] ),
        .I2(\f_permutation_l_/out_reg_n_0_[302] ),
        .I3(\out[1265]_i_2_n_0 ),
        .I4(\out[896]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [704]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[705]_i_1 
       (.I0(\out[1415]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[377] ),
        .I2(\f_permutation_l_/out_reg_n_0_[303] ),
        .I3(\out[1266]_i_2_n_0 ),
        .I4(\out[897]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [705]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[706]_i_1 
       (.I0(\out[1416]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[378] ),
        .I2(\f_permutation_l_/out_reg_n_0_[304] ),
        .I3(\out[1267]_i_2_n_0 ),
        .I4(\out[898]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [706]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[707]_i_1 
       (.I0(\out[1417]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[379] ),
        .I2(\f_permutation_l_/out_reg_n_0_[305] ),
        .I3(\out[1268]_i_2_n_0 ),
        .I4(\out[899]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [707]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[708]_i_1 
       (.I0(\out[1418]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[380] ),
        .I2(\f_permutation_l_/out_reg_n_0_[306] ),
        .I3(\out[1269]_i_2_n_0 ),
        .I4(\out[900]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [708]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[709]_i_1 
       (.I0(\out[1419]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[381] ),
        .I2(\f_permutation_l_/out_reg_n_0_[307] ),
        .I3(\out[1270]_i_2_n_0 ),
        .I4(\out[901]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [709]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[70]_i_1 
       (.I0(\out[1248]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[605] ),
        .I2(\f_permutation_l_/out_reg_n_0_[196] ),
        .I3(\out[1584]_i_3_n_0 ),
        .I4(\out[262]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [70]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[710]_i_1 
       (.I0(\out[1420]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[382] ),
        .I2(\f_permutation_l_/out_reg_n_0_[308] ),
        .I3(\out[1271]_i_2_n_0 ),
        .I4(\out[902]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [710]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[711]_i_1 
       (.I0(\out[1421]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[383] ),
        .I2(\f_permutation_l_/out_reg_n_0_[309] ),
        .I3(\out[1272]_i_2_n_0 ),
        .I4(\out[903]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [711]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[712]_i_1 
       (.I0(\out[1422]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[320] ),
        .I2(\f_permutation_l_/out_reg_n_0_[310] ),
        .I3(\out[1273]_i_2_n_0 ),
        .I4(\out[904]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [712]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[713]_i_1 
       (.I0(\out[1423]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[321] ),
        .I2(\f_permutation_l_/out_reg_n_0_[311] ),
        .I3(\out[1274]_i_2_n_0 ),
        .I4(\out[905]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [713]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[714]_i_1 
       (.I0(\out[1424]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[322] ),
        .I2(\f_permutation_l_/out_reg_n_0_[312] ),
        .I3(\out[1275]_i_2_n_0 ),
        .I4(\out[906]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [714]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[715]_i_1 
       (.I0(\out[1425]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[323] ),
        .I2(\f_permutation_l_/out_reg_n_0_[313] ),
        .I3(\out[1276]_i_2_n_0 ),
        .I4(\out[907]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [715]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[716]_i_1 
       (.I0(\out[1426]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[324] ),
        .I2(\f_permutation_l_/out_reg_n_0_[314] ),
        .I3(\out[1277]_i_2_n_0 ),
        .I4(\out[908]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [716]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[717]_i_1 
       (.I0(\out[1427]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[325] ),
        .I2(\f_permutation_l_/out_reg_n_0_[315] ),
        .I3(\out[1278]_i_2_n_0 ),
        .I4(\out[909]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [717]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[718]_i_1 
       (.I0(\out[1428]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[326] ),
        .I2(\f_permutation_l_/out_reg_n_0_[316] ),
        .I3(\out[1279]_i_2_n_0 ),
        .I4(\out[910]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [718]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[719]_i_1 
       (.I0(\out[1429]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[327] ),
        .I2(\f_permutation_l_/out_reg_n_0_[317] ),
        .I3(\out[1216]_i_2_n_0 ),
        .I4(\out[911]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [719]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[71]_i_1 
       (.I0(\out[1249]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[606] ),
        .I2(\f_permutation_l_/out_reg_n_0_[197] ),
        .I3(\out[1585]_i_3_n_0 ),
        .I4(\out[263]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [71]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[720]_i_1 
       (.I0(\out[1430]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[328] ),
        .I2(\f_permutation_l_/out_reg_n_0_[318] ),
        .I3(\out[1217]_i_2_n_0 ),
        .I4(\out[912]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [720]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[721]_i_1 
       (.I0(\out[1431]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[329] ),
        .I2(\f_permutation_l_/out_reg_n_0_[319] ),
        .I3(\out[1218]_i_2_n_0 ),
        .I4(\out[913]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [721]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[722]_i_1 
       (.I0(\out[1432]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[330] ),
        .I2(\f_permutation_l_/out_reg_n_0_[256] ),
        .I3(\out[1219]_i_2_n_0 ),
        .I4(\out[914]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [722]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[723]_i_1 
       (.I0(\out[1433]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[331] ),
        .I2(\f_permutation_l_/out_reg_n_0_[257] ),
        .I3(\out[1220]_i_2_n_0 ),
        .I4(\out[915]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [723]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[724]_i_1 
       (.I0(\out[1434]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[332] ),
        .I2(\f_permutation_l_/out_reg_n_0_[258] ),
        .I3(\out[1221]_i_2_n_0 ),
        .I4(\out[916]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [724]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[725]_i_1 
       (.I0(\out[1435]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[333] ),
        .I2(\f_permutation_l_/out_reg_n_0_[259] ),
        .I3(\out[1539]_i_6_n_0 ),
        .I4(\out[917]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [725]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[726]_i_1 
       (.I0(\out[1436]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[334] ),
        .I2(\f_permutation_l_/out_reg_n_0_[260] ),
        .I3(\out[1223]_i_2_n_0 ),
        .I4(\out[918]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [726]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[727]_i_1 
       (.I0(\out[1437]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[335] ),
        .I2(\f_permutation_l_/out_reg_n_0_[261] ),
        .I3(\out[1224]_i_2_n_0 ),
        .I4(\out[919]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [727]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[728]_i_1 
       (.I0(\out[1438]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[336] ),
        .I2(\f_permutation_l_/out_reg_n_0_[262] ),
        .I3(\out[1225]_i_2_n_0 ),
        .I4(\out[920]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [728]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[729]_i_1 
       (.I0(\out[1439]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[337] ),
        .I2(\f_permutation_l_/out_reg_n_0_[263] ),
        .I3(\out[1226]_i_2_n_0 ),
        .I4(\out[921]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [729]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[72]_i_1 
       (.I0(\out[1250]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[607] ),
        .I2(\f_permutation_l_/out_reg_n_0_[198] ),
        .I3(\out[1586]_i_3_n_0 ),
        .I4(\out[264]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [72]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[730]_i_1 
       (.I0(\out[1440]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[338] ),
        .I2(\f_permutation_l_/out_reg_n_0_[264] ),
        .I3(\out[1227]_i_2_n_0 ),
        .I4(\out[922]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [730]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[731]_i_1 
       (.I0(\out[1441]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[339] ),
        .I2(\f_permutation_l_/out_reg_n_0_[265] ),
        .I3(\out[1228]_i_2_n_0 ),
        .I4(\out[923]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [731]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[732]_i_1 
       (.I0(\out[1442]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[340] ),
        .I2(\f_permutation_l_/out_reg_n_0_[266] ),
        .I3(\out[1229]_i_2_n_0 ),
        .I4(\out[924]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [732]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[733]_i_1 
       (.I0(\out[1443]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[341] ),
        .I2(\f_permutation_l_/out_reg_n_0_[267] ),
        .I3(\out[1230]_i_2_n_0 ),
        .I4(\out[925]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [733]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[734]_i_1 
       (.I0(\out[1444]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[342] ),
        .I2(\f_permutation_l_/out_reg_n_0_[268] ),
        .I3(\out[1231]_i_2_n_0 ),
        .I4(\out[734]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [734]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[734]_i_2 
       (.I0(\f_permutation_l_/round_in [1501]),
        .I1(\f_permutation_l_/round_in [1436]),
        .I2(\out[1545]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1565]),
        .I4(\out[1545]_i_6_n_0 ),
        .O(\out[734]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[735]_i_1 
       (.I0(\out[1445]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[343] ),
        .I2(\f_permutation_l_/out_reg_n_0_[269] ),
        .I3(\out[1232]_i_2_n_0 ),
        .I4(\out[927]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [735]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[736]_i_1 
       (.I0(\out[1446]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[344] ),
        .I2(\f_permutation_l_/out_reg_n_0_[270] ),
        .I3(\out[1233]_i_2_n_0 ),
        .I4(\out[928]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [736]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[737]_i_1 
       (.I0(\out[1447]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[345] ),
        .I2(\f_permutation_l_/out_reg_n_0_[271] ),
        .I3(\out[1234]_i_2_n_0 ),
        .I4(\out[929]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [737]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[738]_i_1 
       (.I0(\out[1448]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[346] ),
        .I2(\f_permutation_l_/out_reg_n_0_[272] ),
        .I3(\out[1235]_i_2_n_0 ),
        .I4(\out[930]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [738]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[739]_i_1 
       (.I0(\out[1449]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[347] ),
        .I2(\f_permutation_l_/out_reg_n_0_[273] ),
        .I3(\out[1236]_i_2_n_0 ),
        .I4(\out[931]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [739]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[73]_i_1 
       (.I0(\out[1251]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[608] ),
        .I2(\f_permutation_l_/out_reg_n_0_[199] ),
        .I3(\out[1587]_i_3_n_0 ),
        .I4(\out[265]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [73]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[740]_i_1 
       (.I0(\out[1450]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[348] ),
        .I2(\f_permutation_l_/out_reg_n_0_[274] ),
        .I3(\out[1237]_i_2_n_0 ),
        .I4(\out[932]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [740]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[741]_i_1 
       (.I0(\out[1451]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[349] ),
        .I2(\f_permutation_l_/out_reg_n_0_[275] ),
        .I3(\out[1238]_i_2_n_0 ),
        .I4(\out[933]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [741]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[742]_i_1 
       (.I0(\out[1452]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[350] ),
        .I2(\f_permutation_l_/out_reg_n_0_[276] ),
        .I3(\out[1239]_i_2_n_0 ),
        .I4(\out[934]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [742]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[743]_i_1 
       (.I0(\out[1453]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[351] ),
        .I2(\f_permutation_l_/out_reg_n_0_[277] ),
        .I3(\out[1240]_i_2_n_0 ),
        .I4(\out[935]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [743]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696666)) 
    \out[744]_i_1 
       (.I0(\out[1454]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[352] ),
        .I2(\f_permutation_l_/out_reg_n_0_[278] ),
        .I3(\out[1241]_i_2_n_0 ),
        .I4(\out[936]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [744]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[745]_i_1 
       (.I0(\out[1455]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[353] ),
        .I2(\f_permutation_l_/out_reg_n_0_[279] ),
        .I3(\out[1242]_i_2_n_0 ),
        .I4(\out[937]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [745]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[746]_i_1 
       (.I0(\out[1456]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[354] ),
        .I2(\f_permutation_l_/out_reg_n_0_[280] ),
        .I3(\out[1243]_i_2_n_0 ),
        .I4(\out[938]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [746]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[747]_i_1 
       (.I0(\out[1457]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[355] ),
        .I2(\f_permutation_l_/out_reg_n_0_[281] ),
        .I3(\out[1244]_i_2_n_0 ),
        .I4(\out[939]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [747]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[748]_i_1 
       (.I0(\out[1458]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[356] ),
        .I2(\f_permutation_l_/out_reg_n_0_[282] ),
        .I3(\out[1245]_i_2_n_0 ),
        .I4(\out[940]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [748]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[749]_i_1 
       (.I0(\out[1459]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[357] ),
        .I2(\f_permutation_l_/out_reg_n_0_[283] ),
        .I3(\out[1246]_i_2_n_0 ),
        .I4(\out[941]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [749]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[74]_i_1 
       (.I0(\out[1252]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[609] ),
        .I2(\f_permutation_l_/out_reg_n_0_[200] ),
        .I3(\out[1588]_i_3_n_0 ),
        .I4(\out[266]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [74]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[750]_i_1 
       (.I0(\out[1460]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[358] ),
        .I2(\f_permutation_l_/out_reg_n_0_[284] ),
        .I3(\out[1247]_i_2_n_0 ),
        .I4(\out[942]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [750]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[751]_i_1 
       (.I0(\out[1461]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[359] ),
        .I2(\f_permutation_l_/out_reg_n_0_[285] ),
        .I3(\out[1248]_i_2_n_0 ),
        .I4(\out[943]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [751]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[752]_i_1 
       (.I0(\out[1462]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[360] ),
        .I2(\f_permutation_l_/out_reg_n_0_[286] ),
        .I3(\out[1249]_i_2_n_0 ),
        .I4(\out[944]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [752]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[753]_i_1 
       (.I0(\out[1463]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[361] ),
        .I2(\f_permutation_l_/out_reg_n_0_[287] ),
        .I3(\out[1250]_i_2_n_0 ),
        .I4(\out[945]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [753]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[754]_i_1 
       (.I0(\out[1464]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[362] ),
        .I2(\f_permutation_l_/out_reg_n_0_[288] ),
        .I3(\out[1251]_i_2_n_0 ),
        .I4(\out[946]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [754]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[755]_i_1 
       (.I0(\out[1465]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[363] ),
        .I2(\f_permutation_l_/out_reg_n_0_[289] ),
        .I3(\out[1252]_i_2_n_0 ),
        .I4(\out[947]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [755]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[756]_i_1 
       (.I0(\out[1466]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[364] ),
        .I2(\f_permutation_l_/out_reg_n_0_[290] ),
        .I3(\out[1253]_i_2_n_0 ),
        .I4(\out[948]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [756]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[757]_i_1 
       (.I0(\out[1467]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[365] ),
        .I2(\f_permutation_l_/out_reg_n_0_[291] ),
        .I3(\out[1254]_i_2_n_0 ),
        .I4(\out[949]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [757]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[758]_i_1 
       (.I0(\out[1468]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[366] ),
        .I2(\f_permutation_l_/out_reg_n_0_[292] ),
        .I3(\out[1255]_i_2_n_0 ),
        .I4(\out[950]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [758]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[759]_i_1 
       (.I0(\out[1469]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[367] ),
        .I2(\f_permutation_l_/out_reg_n_0_[293] ),
        .I3(\out[1256]_i_2_n_0 ),
        .I4(\out[951]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [759]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[75]_i_1 
       (.I0(\out[1253]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[610] ),
        .I2(\f_permutation_l_/out_reg_n_0_[201] ),
        .I3(\out[1589]_i_3_n_0 ),
        .I4(\out[267]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [75]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[760]_i_1 
       (.I0(\out[1470]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[368] ),
        .I2(\f_permutation_l_/out_reg_n_0_[294] ),
        .I3(\out[1257]_i_2_n_0 ),
        .I4(\out[952]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [760]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[761]_i_1 
       (.I0(\out[1471]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[369] ),
        .I2(\f_permutation_l_/out_reg_n_0_[295] ),
        .I3(\out[1258]_i_2_n_0 ),
        .I4(\out[953]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [761]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[762]_i_1 
       (.I0(\out[1408]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[370] ),
        .I2(\f_permutation_l_/out_reg_n_0_[296] ),
        .I3(\out[1259]_i_2_n_0 ),
        .I4(\out[954]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [762]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[763]_i_1 
       (.I0(\out[1409]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[371] ),
        .I2(\f_permutation_l_/out_reg_n_0_[297] ),
        .I3(\out[1260]_i_2_n_0 ),
        .I4(\out[955]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [763]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[764]_i_1 
       (.I0(\out[1410]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[372] ),
        .I2(\f_permutation_l_/out_reg_n_0_[298] ),
        .I3(\out[1261]_i_2_n_0 ),
        .I4(\out[956]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [764]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[765]_i_1 
       (.I0(\out[1411]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[373] ),
        .I2(\f_permutation_l_/out_reg_n_0_[299] ),
        .I3(\out[1262]_i_2_n_0 ),
        .I4(\out[957]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [765]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[766]_i_1 
       (.I0(\out[1412]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[374] ),
        .I2(\f_permutation_l_/out_reg_n_0_[300] ),
        .I3(\out[1263]_i_2_n_0 ),
        .I4(\out[958]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [766]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69966666)) 
    \out[767]_i_1 
       (.I0(\out[1413]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[375] ),
        .I2(\f_permutation_l_/out_reg_n_0_[301] ),
        .I3(\out[1264]_i_2_n_0 ),
        .I4(\out[959]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [767]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[768]_i_1 
       (.I0(\out[1532]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[743] ),
        .I2(\out[768]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[302] ),
        .I4(\out[1265]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [768]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[768]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[376] ),
        .I1(\out[1571]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1591]),
        .I3(\f_permutation_l_/round_in [1400]),
        .I4(\out[1572]_i_10_n_0 ),
        .O(\out[768]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[769]_i_1 
       (.I0(\out[1533]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[744] ),
        .I2(\out[769]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[303] ),
        .I4(\out[1266]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [769]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[769]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[377] ),
        .I1(\out[1572]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1592]),
        .I3(\f_permutation_l_/round_in [1401]),
        .I4(\out[1573]_i_10_n_0 ),
        .O(\out[769]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[76]_i_1 
       (.I0(\out[1254]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[611] ),
        .I2(\f_permutation_l_/out_reg_n_0_[202] ),
        .I3(\out[1590]_i_3_n_0 ),
        .I4(\out[268]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [76]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[770]_i_1 
       (.I0(\out[1534]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[745] ),
        .I2(\out[770]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[304] ),
        .I4(\out[1267]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [770]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[770]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[378] ),
        .I1(\out[1573]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1593]),
        .I3(\f_permutation_l_/round_in [1402]),
        .I4(\out[1574]_i_10_n_0 ),
        .O(\out[770]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[771]_i_1 
       (.I0(\out[1535]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[746] ),
        .I2(\out[771]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[305] ),
        .I4(\out[1268]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [771]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[771]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[379] ),
        .I1(\out[1574]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1594]),
        .I3(\f_permutation_l_/round_in [1403]),
        .I4(\out[1575]_i_10_n_0 ),
        .O(\out[771]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[772]_i_1 
       (.I0(\out[1472]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[747] ),
        .I2(\out[772]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[306] ),
        .I4(\out[1269]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [772]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[772]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[380] ),
        .I1(\out[1575]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1595]),
        .I3(\f_permutation_l_/round_in [1404]),
        .I4(\out[1576]_i_10_n_0 ),
        .O(\out[772]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[773]_i_1 
       (.I0(\out[1473]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[748] ),
        .I2(\out[773]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[307] ),
        .I4(\out[1270]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [773]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[773]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[381] ),
        .I1(\out[1576]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1596]),
        .I3(\f_permutation_l_/round_in [1405]),
        .I4(\out[1577]_i_10_n_0 ),
        .O(\out[773]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[774]_i_1 
       (.I0(\out[1474]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[749] ),
        .I2(\out[774]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[308] ),
        .I4(\out[1271]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [774]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[774]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[382] ),
        .I1(\f_permutation_l_/round_in [1597]),
        .I2(\out[1577]_i_6_n_0 ),
        .I3(\out[1578]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1406]),
        .O(\out[774]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[775]_i_1 
       (.I0(\out[1475]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[750] ),
        .I2(\out[775]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[309] ),
        .I4(\out[1272]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [775]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[775]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[383] ),
        .I1(\f_permutation_l_/round_in [1598]),
        .I2(\out[1578]_i_6_n_0 ),
        .I3(\out[1579]_i_10_n_0 ),
        .I4(\f_permutation_l_/round_in [1407]),
        .O(\out[775]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[776]_i_1 
       (.I0(\out[1476]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[751] ),
        .I2(\out[776]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[310] ),
        .I4(\out[1273]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [776]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[776]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[320] ),
        .I1(\f_permutation_l_/round_in [1599]),
        .I2(\out[1579]_i_7_n_0 ),
        .I3(\out[1580]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1344]),
        .O(\out[776]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[777]_i_1 
       (.I0(\out[1477]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[752] ),
        .I2(\out[777]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[311] ),
        .I4(\out[1274]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [777]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[777]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[321] ),
        .I1(\f_permutation_l_/round_in [1536]),
        .I2(\out[1580]_i_6_n_0 ),
        .I3(\out[1581]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1345]),
        .O(\out[777]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[778]_i_1 
       (.I0(\out[1478]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[753] ),
        .I2(\out[778]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[312] ),
        .I4(\out[1275]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [778]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[778]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[322] ),
        .I1(\f_permutation_l_/round_in [1537]),
        .I2(\out[1581]_i_6_n_0 ),
        .I3(\out[1582]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1346]),
        .O(\out[778]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[779]_i_1 
       (.I0(\out[1479]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[754] ),
        .I2(\out[779]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[313] ),
        .I4(\out[1276]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [779]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[779]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[323] ),
        .I1(\f_permutation_l_/round_in [1538]),
        .I2(\out[1582]_i_6_n_0 ),
        .I3(\out[1583]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1347]),
        .O(\out[779]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[77]_i_1 
       (.I0(\out[1255]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[612] ),
        .I2(\f_permutation_l_/out_reg_n_0_[203] ),
        .I3(\out[1591]_i_3_n_0 ),
        .I4(\out[269]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [77]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[780]_i_1 
       (.I0(\out[1480]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[755] ),
        .I2(\out[780]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[314] ),
        .I4(\out[1277]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [780]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[780]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[324] ),
        .I1(\f_permutation_l_/round_in [1539]),
        .I2(\out[1583]_i_6_n_0 ),
        .I3(\out[1584]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1348]),
        .O(\out[780]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[781]_i_1 
       (.I0(\out[1481]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[756] ),
        .I2(\out[781]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[315] ),
        .I4(\out[1278]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [781]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[781]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[325] ),
        .I1(\f_permutation_l_/round_in [1540]),
        .I2(\out[1584]_i_6_n_0 ),
        .I3(\out[1585]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1349]),
        .O(\out[781]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[782]_i_1 
       (.I0(\out[1482]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[757] ),
        .I2(\out[782]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[316] ),
        .I4(\out[1279]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [782]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[782]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[326] ),
        .I1(\f_permutation_l_/round_in [1541]),
        .I2(\out[1585]_i_6_n_0 ),
        .I3(\out[1586]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1350]),
        .O(\out[782]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[783]_i_1 
       (.I0(\out[1483]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[758] ),
        .I2(\out[783]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[317] ),
        .I4(\out[1216]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [783]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[783]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[327] ),
        .I1(\f_permutation_l_/round_in [1542]),
        .I2(\out[1586]_i_6_n_0 ),
        .I3(\out[1587]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1351]),
        .O(\out[783]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[784]_i_1 
       (.I0(\out[1484]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[759] ),
        .I2(\out[784]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[318] ),
        .I4(\out[1217]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [784]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[784]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[328] ),
        .I1(\f_permutation_l_/round_in [1543]),
        .I2(\out[1587]_i_6_n_0 ),
        .I3(\out[1588]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1352]),
        .O(\out[784]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[785]_i_1 
       (.I0(\out[1485]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[760] ),
        .I2(\out[785]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[319] ),
        .I4(\out[1218]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [785]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[785]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[329] ),
        .I1(\f_permutation_l_/round_in [1544]),
        .I2(\out[1588]_i_6_n_0 ),
        .I3(\out[1589]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1353]),
        .O(\out[785]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[786]_i_1 
       (.I0(\out[1486]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[761] ),
        .I2(\out[786]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[256] ),
        .I4(\out[1219]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [786]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[786]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[330] ),
        .I1(\f_permutation_l_/round_in [1545]),
        .I2(\out[1589]_i_6_n_0 ),
        .I3(\out[1590]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1354]),
        .O(\out[786]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[787]_i_1 
       (.I0(\out[1487]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[762] ),
        .I2(\out[787]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[257] ),
        .I4(\out[1220]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [787]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[787]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[331] ),
        .I1(\f_permutation_l_/round_in [1546]),
        .I2(\out[1590]_i_6_n_0 ),
        .I3(\out[1591]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1355]),
        .O(\out[787]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[788]_i_1 
       (.I0(\out[1488]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[763] ),
        .I2(\out[788]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[258] ),
        .I4(\out[1221]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [788]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[788]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[332] ),
        .I1(\f_permutation_l_/round_in [1547]),
        .I2(\out[1591]_i_6_n_0 ),
        .I3(\out[1592]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1356]),
        .O(\out[788]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[789]_i_1 
       (.I0(\out[1489]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[764] ),
        .I2(\out[789]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[259] ),
        .I4(\out[1539]_i_6_n_0 ),
        .O(\f_permutation_l_/round_out [789]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[789]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[333] ),
        .I1(\f_permutation_l_/round_in [1548]),
        .I2(\out[1592]_i_6_n_0 ),
        .I3(\out[1593]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1357]),
        .O(\out[789]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[78]_i_1 
       (.I0(\out[1256]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[613] ),
        .I2(\f_permutation_l_/out_reg_n_0_[204] ),
        .I3(\out[1592]_i_3_n_0 ),
        .I4(\out[270]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [78]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[790]_i_1 
       (.I0(\out[1490]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[765] ),
        .I2(\out[790]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[260] ),
        .I4(\out[1223]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [790]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[790]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[334] ),
        .I1(\f_permutation_l_/round_in [1549]),
        .I2(\out[1593]_i_6_n_0 ),
        .I3(\out[1594]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1358]),
        .O(\out[790]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[791]_i_1 
       (.I0(\out[1491]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[766] ),
        .I2(\out[791]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[261] ),
        .I4(\out[1224]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [791]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[791]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[335] ),
        .I1(\f_permutation_l_/round_in [1550]),
        .I2(\out[1594]_i_6_n_0 ),
        .I3(\out[1595]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1359]),
        .O(\out[791]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[792]_i_1 
       (.I0(\out[1492]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[767] ),
        .I2(\out[792]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[262] ),
        .I4(\out[1225]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [792]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[792]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[336] ),
        .I1(\f_permutation_l_/round_in [1551]),
        .I2(\out[1595]_i_6_n_0 ),
        .I3(\out[1596]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1360]),
        .O(\out[792]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[793]_i_1 
       (.I0(\out[1493]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[704] ),
        .I2(\out[793]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[263] ),
        .I4(\out[1226]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [793]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[793]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[337] ),
        .I1(\f_permutation_l_/round_in [1552]),
        .I2(\out[1596]_i_6_n_0 ),
        .I3(\out[1597]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1361]),
        .O(\out[793]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[794]_i_1 
       (.I0(\out[1494]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[705] ),
        .I2(\out[794]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[264] ),
        .I4(\out[1227]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [794]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[794]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[338] ),
        .I1(\f_permutation_l_/round_in [1553]),
        .I2(\out[1597]_i_6_n_0 ),
        .I3(\out[1598]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1362]),
        .O(\out[794]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[795]_i_1 
       (.I0(\out[1495]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[706] ),
        .I2(\out[795]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[265] ),
        .I4(\out[1228]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [795]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[795]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[339] ),
        .I1(\f_permutation_l_/round_in [1554]),
        .I2(\out[1598]_i_6_n_0 ),
        .I3(\out[1599]_i_9_n_0 ),
        .I4(\f_permutation_l_/round_in [1363]),
        .O(\out[795]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[796]_i_1 
       (.I0(\out[1496]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[707] ),
        .I2(\out[796]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[266] ),
        .I4(\out[1229]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [796]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[796]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[340] ),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1555]),
        .I4(\out[1599]_i_8_n_0 ),
        .O(\out[796]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[797]_i_1 
       (.I0(\out[1497]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[708] ),
        .I2(\out[797]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[267] ),
        .I4(\out[1230]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [797]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[797]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[341] ),
        .I1(\out[1536]_i_10_n_0 ),
        .I2(\f_permutation_l_/round_in [1556]),
        .I3(\f_permutation_l_/round_in [1365]),
        .I4(\out[1537]_i_11_n_0 ),
        .O(\out[797]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[798]_i_1 
       (.I0(\out[1498]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[709] ),
        .I2(\out[798]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[268] ),
        .I4(\out[1231]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [798]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[798]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[342] ),
        .I1(\out[1537]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1557]),
        .I3(\f_permutation_l_/round_in [1366]),
        .I4(\out[1538]_i_10_n_0 ),
        .O(\out[798]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[799]_i_1 
       (.I0(\out[1499]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[710] ),
        .I2(\out[799]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[269] ),
        .I4(\out[1232]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [799]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[799]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[343] ),
        .I1(\f_permutation_l_/round_in [1558]),
        .I2(\out[1538]_i_6_n_0 ),
        .I3(\out[1539]_i_12_n_0 ),
        .I4(\f_permutation_l_/round_in [1367]),
        .O(\out[799]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[79]_i_1 
       (.I0(\out[1257]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[614] ),
        .I2(\f_permutation_l_/out_reg_n_0_[205] ),
        .I3(\out[1593]_i_3_n_0 ),
        .I4(\out[271]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [79]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[7]_i_1 
       (.I0(\out[1585]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[197] ),
        .I2(\out[263]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1040]),
        .I4(\out[1509]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[800]_i_1 
       (.I0(\out[1500]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[711] ),
        .I2(\out[800]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[270] ),
        .I4(\out[1233]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [800]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[800]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[344] ),
        .I1(\out[1539]_i_8_n_0 ),
        .I2(\f_permutation_l_/round_in [1559]),
        .I3(\f_permutation_l_/round_in [1368]),
        .I4(\out[1540]_i_10_n_0 ),
        .O(\out[800]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[801]_i_1 
       (.I0(\out[1501]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[712] ),
        .I2(\out[801]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[271] ),
        .I4(\out[1234]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [801]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[801]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[345] ),
        .I1(\out[1540]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1560]),
        .I3(\f_permutation_l_/round_in [1369]),
        .I4(\out[1541]_i_10_n_0 ),
        .O(\out[801]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[802]_i_1 
       (.I0(\out[1502]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[713] ),
        .I2(\out[802]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[272] ),
        .I4(\out[1235]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [802]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[802]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[346] ),
        .I1(\out[1541]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1561]),
        .I3(\f_permutation_l_/round_in [1370]),
        .I4(\out[1542]_i_12_n_0 ),
        .O(\out[802]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[803]_i_1 
       (.I0(\out[1503]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[714] ),
        .I2(\out[803]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[273] ),
        .I4(\out[1236]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [803]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[803]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[347] ),
        .I1(\out[1542]_i_7_n_0 ),
        .I2(\f_permutation_l_/round_in [1562]),
        .I3(\f_permutation_l_/round_in [1371]),
        .I4(\out[1543]_i_13_n_0 ),
        .O(\out[803]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[804]_i_1 
       (.I0(\out[1504]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[715] ),
        .I2(\out[804]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[274] ),
        .I4(\out[1237]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [804]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[804]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[348] ),
        .I1(\out[1543]_i_10_n_0 ),
        .I2(\f_permutation_l_/round_in [1563]),
        .I3(\f_permutation_l_/round_in [1372]),
        .I4(\out[1544]_i_10_n_0 ),
        .O(\out[804]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[805]_i_1 
       (.I0(\out[1505]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[716] ),
        .I2(\out[805]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[275] ),
        .I4(\out[1238]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [805]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[805]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[349] ),
        .I1(\out[1544]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1564]),
        .I3(\f_permutation_l_/round_in [1373]),
        .I4(\out[1545]_i_10_n_0 ),
        .O(\out[805]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[806]_i_1 
       (.I0(\out[1506]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[717] ),
        .I2(\out[806]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[276] ),
        .I4(\out[1239]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [806]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[806]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[350] ),
        .I1(\out[1545]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1565]),
        .I3(\f_permutation_l_/round_in [1374]),
        .I4(\out[1546]_i_10_n_0 ),
        .O(\out[806]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[807]_i_1 
       (.I0(\out[1507]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[718] ),
        .I2(\out[807]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[277] ),
        .I4(\out[1240]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [807]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[807]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[351] ),
        .I1(\out[1546]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1566]),
        .I3(\f_permutation_l_/round_in [1375]),
        .I4(\out[1547]_i_10_n_0 ),
        .O(\out[807]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[808]_i_1 
       (.I0(\out[1508]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[719] ),
        .I2(\out[808]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[278] ),
        .I4(\out[1241]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [808]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[808]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[352] ),
        .I1(\out[1547]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1567]),
        .I3(\f_permutation_l_/round_in [1376]),
        .I4(\out[1548]_i_10_n_0 ),
        .O(\out[808]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[809]_i_1 
       (.I0(\out[1509]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[720] ),
        .I2(\out[809]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[279] ),
        .I4(\out[1242]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [809]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[809]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[353] ),
        .I1(\out[1548]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1568]),
        .I3(\f_permutation_l_/round_in [1377]),
        .I4(\out[1549]_i_10_n_0 ),
        .O(\out[809]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[80]_i_1 
       (.I0(\out[1258]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[615] ),
        .I2(\f_permutation_l_/out_reg_n_0_[206] ),
        .I3(\out[1594]_i_3_n_0 ),
        .I4(\out[272]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [80]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[810]_i_1 
       (.I0(\out[1510]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[721] ),
        .I2(\out[810]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[280] ),
        .I4(\out[1243]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [810]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[810]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[354] ),
        .I1(\out[1549]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1569]),
        .I3(\f_permutation_l_/round_in [1378]),
        .I4(\out[1550]_i_10_n_0 ),
        .O(\out[810]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[811]_i_1 
       (.I0(\out[1511]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[722] ),
        .I2(\out[811]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[281] ),
        .I4(\out[1244]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [811]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[811]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[355] ),
        .I1(\out[1550]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1570]),
        .I3(\f_permutation_l_/round_in [1379]),
        .I4(\out[1551]_i_11_n_0 ),
        .O(\out[811]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[812]_i_1 
       (.I0(\out[1512]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[723] ),
        .I2(\out[812]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[282] ),
        .I4(\out[1245]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [812]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[812]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[356] ),
        .I1(\out[1551]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1571]),
        .I3(\f_permutation_l_/round_in [1380]),
        .I4(\out[1552]_i_10_n_0 ),
        .O(\out[812]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[813]_i_1 
       (.I0(\out[1513]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[724] ),
        .I2(\out[813]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[283] ),
        .I4(\out[1246]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [813]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[813]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[357] ),
        .I1(\out[1552]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1572]),
        .I3(\f_permutation_l_/round_in [1381]),
        .I4(\out[1553]_i_10_n_0 ),
        .O(\out[813]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[814]_i_1 
       (.I0(\out[1514]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[725] ),
        .I2(\out[814]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[284] ),
        .I4(\out[1247]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [814]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[814]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[358] ),
        .I1(\out[1553]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1573]),
        .I3(\f_permutation_l_/round_in [1382]),
        .I4(\out[1554]_i_10_n_0 ),
        .O(\out[814]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69666669)) 
    \out[815]_i_1 
       (.I0(\out[1515]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[726] ),
        .I2(\out[815]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[285] ),
        .I4(\out[1248]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [815]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[815]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[359] ),
        .I1(\out[1554]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1574]),
        .I3(\f_permutation_l_/round_in [1383]),
        .I4(\out[1555]_i_10_n_0 ),
        .O(\out[815]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[816]_i_1 
       (.I0(\out[1516]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[727] ),
        .I2(\out[816]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[286] ),
        .I4(\out[1249]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [816]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[816]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[360] ),
        .I1(\out[1555]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1575]),
        .I3(\f_permutation_l_/round_in [1384]),
        .I4(\out[1556]_i_11_n_0 ),
        .O(\out[816]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[817]_i_1 
       (.I0(\out[1517]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[728] ),
        .I2(\out[817]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[287] ),
        .I4(\out[1250]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [817]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[817]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[361] ),
        .I1(\out[1556]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1576]),
        .I3(\f_permutation_l_/round_in [1385]),
        .I4(\out[1557]_i_10_n_0 ),
        .O(\out[817]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[818]_i_1 
       (.I0(\out[1518]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[729] ),
        .I2(\out[818]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[288] ),
        .I4(\out[1251]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [818]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[818]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[362] ),
        .I1(\out[1557]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1577]),
        .I3(\f_permutation_l_/round_in [1386]),
        .I4(\out[1558]_i_10_n_0 ),
        .O(\out[818]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[819]_i_1 
       (.I0(\out[1519]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[730] ),
        .I2(\out[819]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[289] ),
        .I4(\out[1252]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [819]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[819]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[363] ),
        .I1(\out[1558]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1578]),
        .I3(\f_permutation_l_/round_in [1387]),
        .I4(\out[1559]_i_10_n_0 ),
        .O(\out[819]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[81]_i_1 
       (.I0(\out[1259]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[616] ),
        .I2(\f_permutation_l_/out_reg_n_0_[207] ),
        .I3(\out[1595]_i_3_n_0 ),
        .I4(\out[273]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [81]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[820]_i_1 
       (.I0(\out[1520]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[731] ),
        .I2(\out[820]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[290] ),
        .I4(\out[1253]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [820]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[820]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[364] ),
        .I1(\out[1559]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1579]),
        .I3(\f_permutation_l_/round_in [1388]),
        .I4(\out[1560]_i_10_n_0 ),
        .O(\out[820]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[821]_i_1 
       (.I0(\out[1521]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[732] ),
        .I2(\out[821]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[291] ),
        .I4(\out[1254]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [821]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[821]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[365] ),
        .I1(\out[1560]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1580]),
        .I3(\f_permutation_l_/round_in [1389]),
        .I4(\out[1561]_i_10_n_0 ),
        .O(\out[821]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[822]_i_1 
       (.I0(\out[1522]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[733] ),
        .I2(\out[822]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[292] ),
        .I4(\out[1255]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [822]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[822]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[366] ),
        .I1(\out[1561]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1581]),
        .I3(\f_permutation_l_/round_in [1390]),
        .I4(\out[1562]_i_10_n_0 ),
        .O(\out[822]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[823]_i_1 
       (.I0(\out[1523]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[734] ),
        .I2(\out[823]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[293] ),
        .I4(\out[1256]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [823]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[823]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[367] ),
        .I1(\out[1562]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1582]),
        .I3(\f_permutation_l_/round_in [1391]),
        .I4(\out[1563]_i_10_n_0 ),
        .O(\out[823]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[824]_i_1 
       (.I0(\out[1524]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[735] ),
        .I2(\out[824]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[294] ),
        .I4(\out[1257]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [824]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[824]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[368] ),
        .I1(\out[1563]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1583]),
        .I3(\f_permutation_l_/round_in [1392]),
        .I4(\out[1564]_i_10_n_0 ),
        .O(\out[824]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[825]_i_1 
       (.I0(\out[1525]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[736] ),
        .I2(\out[825]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[295] ),
        .I4(\out[1258]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [825]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[825]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[369] ),
        .I1(\out[1564]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1584]),
        .I3(\f_permutation_l_/round_in [1393]),
        .I4(\out[1565]_i_10_n_0 ),
        .O(\out[825]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[826]_i_1 
       (.I0(\out[1526]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[737] ),
        .I2(\out[826]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[296] ),
        .I4(\out[1259]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [826]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[826]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[370] ),
        .I1(\out[1565]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1585]),
        .I3(\f_permutation_l_/round_in [1394]),
        .I4(\out[1566]_i_10_n_0 ),
        .O(\out[826]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[827]_i_1 
       (.I0(\out[1527]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[738] ),
        .I2(\out[827]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[297] ),
        .I4(\out[1260]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [827]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[827]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[371] ),
        .I1(\out[1566]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1586]),
        .I3(\f_permutation_l_/round_in [1395]),
        .I4(\out[1567]_i_11_n_0 ),
        .O(\out[827]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[828]_i_1 
       (.I0(\out[1528]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[739] ),
        .I2(\out[828]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[298] ),
        .I4(\out[1261]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [828]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[828]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[372] ),
        .I1(\out[1567]_i_9_n_0 ),
        .I2(\f_permutation_l_/round_in [1587]),
        .I3(\f_permutation_l_/round_in [1396]),
        .I4(\out[1568]_i_10_n_0 ),
        .O(\out[828]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[829]_i_1 
       (.I0(\out[1529]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[740] ),
        .I2(\out[829]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[299] ),
        .I4(\out[1262]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [829]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[829]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[373] ),
        .I1(\out[1568]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1588]),
        .I3(\f_permutation_l_/round_in [1397]),
        .I4(\out[1569]_i_10_n_0 ),
        .O(\out[829]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[82]_i_1 
       (.I0(\out[1260]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[617] ),
        .I2(\f_permutation_l_/out_reg_n_0_[208] ),
        .I3(\out[1596]_i_3_n_0 ),
        .I4(\out[274]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [82]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[830]_i_1 
       (.I0(\out[1530]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[741] ),
        .I2(\out[830]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[300] ),
        .I4(\out[1263]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [830]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[830]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[374] ),
        .I1(\out[1569]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1589]),
        .I3(\f_permutation_l_/round_in [1398]),
        .I4(\out[1570]_i_10_n_0 ),
        .O(\out[830]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[831]_i_1 
       (.I0(\out[1531]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[742] ),
        .I2(\out[831]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[301] ),
        .I4(\out[1264]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [831]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[831]_i_2 
       (.I0(\f_permutation_l_/out_reg_n_0_[375] ),
        .I1(\out[1570]_i_6_n_0 ),
        .I2(\f_permutation_l_/round_in [1590]),
        .I3(\f_permutation_l_/round_in [1399]),
        .I4(\out[1571]_i_10_n_0 ),
        .O(\out[831]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[832]_i_1 
       (.I0(\out[832]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[743] ),
        .I2(\out[1532]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[376] ),
        .I4(\out[1414]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [832]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[832]_i_2 
       (.I0(\f_permutation_l_/round_in [1146]),
        .I1(\f_permutation_l_/round_in [1401]),
        .I2(\out[1573]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1530]),
        .I4(\out[1573]_i_9_n_0 ),
        .O(\out[832]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[833]_i_1 
       (.I0(\out[833]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[744] ),
        .I2(\out[1533]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[377] ),
        .I4(\out[1415]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [833]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[833]_i_2 
       (.I0(\f_permutation_l_/round_in [1147]),
        .I1(\f_permutation_l_/round_in [1402]),
        .I2(\out[1574]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1531]),
        .I4(\out[1574]_i_9_n_0 ),
        .O(\out[833]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[834]_i_1 
       (.I0(\out[834]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[745] ),
        .I2(\out[1534]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[378] ),
        .I4(\out[1416]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [834]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[834]_i_2 
       (.I0(\f_permutation_l_/round_in [1148]),
        .I1(\f_permutation_l_/round_in [1403]),
        .I2(\out[1575]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1532]),
        .I4(\out[1575]_i_9_n_0 ),
        .O(\out[834]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[835]_i_1 
       (.I0(\out[835]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[746] ),
        .I2(\out[1535]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[379] ),
        .I4(\out[1417]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [835]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[835]_i_2 
       (.I0(\f_permutation_l_/round_in [1149]),
        .I1(\f_permutation_l_/round_in [1404]),
        .I2(\out[1576]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1533]),
        .I4(\out[1576]_i_9_n_0 ),
        .O(\out[835]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[836]_i_1 
       (.I0(\out[836]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[747] ),
        .I2(\out[1472]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[380] ),
        .I4(\out[1418]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [836]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[836]_i_2 
       (.I0(\f_permutation_l_/round_in [1150]),
        .I1(\f_permutation_l_/round_in [1405]),
        .I2(\out[1577]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1534]),
        .I4(\out[1577]_i_9_n_0 ),
        .O(\out[836]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[837]_i_1 
       (.I0(\out[837]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[748] ),
        .I2(\out[1473]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[381] ),
        .I4(\out[1419]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [837]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[837]_i_2 
       (.I0(\f_permutation_l_/round_in [1151]),
        .I1(\f_permutation_l_/round_in [1406]),
        .I2(\out[1578]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1535]),
        .I4(\out[1536]_i_19_n_0 ),
        .O(\out[837]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[838]_i_1 
       (.I0(\out[838]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[749] ),
        .I2(\out[1474]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[382] ),
        .I4(\out[1420]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [838]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[838]_i_2 
       (.I0(\f_permutation_l_/round_in [1088]),
        .I1(\f_permutation_l_/round_in [1407]),
        .I2(\out[1579]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1472]),
        .I4(\out[1537]_i_17_n_0 ),
        .O(\out[838]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[839]_i_1 
       (.I0(\out[839]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[750] ),
        .I2(\out[1475]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[383] ),
        .I4(\out[1421]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [839]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[839]_i_2 
       (.I0(\f_permutation_l_/round_in [1089]),
        .I1(\f_permutation_l_/round_in [1344]),
        .I2(\out[1580]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1473]),
        .I4(\out[1538]_i_16_n_0 ),
        .O(\out[839]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[83]_i_1 
       (.I0(\out[1261]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[618] ),
        .I2(\f_permutation_l_/out_reg_n_0_[209] ),
        .I3(\out[1597]_i_3_n_0 ),
        .I4(\out[275]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [83]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[840]_i_1 
       (.I0(\out[840]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[751] ),
        .I2(\out[1476]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[320] ),
        .I4(\out[1422]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [840]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[840]_i_2 
       (.I0(\f_permutation_l_/round_in [1090]),
        .I1(\f_permutation_l_/round_in [1345]),
        .I2(\out[1581]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1474]),
        .I4(\out[1539]_i_15_n_0 ),
        .O(\out[840]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[841]_i_1 
       (.I0(\out[841]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[752] ),
        .I2(\out[1477]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[321] ),
        .I4(\out[1423]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [841]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[841]_i_2 
       (.I0(\f_permutation_l_/round_in [1091]),
        .I1(\f_permutation_l_/round_in [1346]),
        .I2(\out[1582]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1475]),
        .I4(\out[1540]_i_16_n_0 ),
        .O(\out[841]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[842]_i_1 
       (.I0(\out[842]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[753] ),
        .I2(\out[1478]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[322] ),
        .I4(\out[1424]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [842]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[842]_i_2 
       (.I0(\f_permutation_l_/round_in [1092]),
        .I1(\f_permutation_l_/round_in [1347]),
        .I2(\out[1583]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1476]),
        .I4(\out[1541]_i_16_n_0 ),
        .O(\out[842]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[843]_i_1 
       (.I0(\out[843]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[754] ),
        .I2(\out[1479]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[323] ),
        .I4(\out[1425]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [843]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[843]_i_2 
       (.I0(\f_permutation_l_/round_in [1093]),
        .I1(\f_permutation_l_/round_in [1348]),
        .I2(\out[1584]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1477]),
        .I4(\out[1542]_i_18_n_0 ),
        .O(\out[843]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[844]_i_1 
       (.I0(\out[844]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[755] ),
        .I2(\out[1480]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[324] ),
        .I4(\out[1426]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [844]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[844]_i_2 
       (.I0(\f_permutation_l_/round_in [1094]),
        .I1(\f_permutation_l_/round_in [1349]),
        .I2(\out[1585]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1478]),
        .I4(\out[1543]_i_19_n_0 ),
        .O(\out[844]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[845]_i_1 
       (.I0(\out[845]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[756] ),
        .I2(\out[1481]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[325] ),
        .I4(\out[1427]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [845]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[845]_i_2 
       (.I0(\f_permutation_l_/round_in [1095]),
        .I1(\f_permutation_l_/round_in [1350]),
        .I2(\out[1586]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1479]),
        .I4(\out[1544]_i_16_n_0 ),
        .O(\out[845]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[846]_i_1 
       (.I0(\out[846]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[757] ),
        .I2(\out[1482]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[326] ),
        .I4(\out[1428]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [846]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[846]_i_2 
       (.I0(\f_permutation_l_/round_in [1096]),
        .I1(\f_permutation_l_/round_in [1351]),
        .I2(\out[1587]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1480]),
        .I4(\out[1545]_i_16_n_0 ),
        .O(\out[846]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[847]_i_1 
       (.I0(\out[847]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[758] ),
        .I2(\out[1483]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[327] ),
        .I4(\out[1429]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [847]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[847]_i_2 
       (.I0(\f_permutation_l_/round_in [1097]),
        .I1(\f_permutation_l_/round_in [1352]),
        .I2(\out[1588]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1481]),
        .I4(\out[1546]_i_16_n_0 ),
        .O(\out[847]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[848]_i_1 
       (.I0(\out[848]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[759] ),
        .I2(\out[1484]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[328] ),
        .I4(\out[1430]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [848]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[848]_i_2 
       (.I0(\f_permutation_l_/round_in [1098]),
        .I1(\f_permutation_l_/round_in [1353]),
        .I2(\out[1589]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1482]),
        .I4(\out[1547]_i_16_n_0 ),
        .O(\out[848]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[849]_i_1 
       (.I0(\out[849]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[760] ),
        .I2(\out[1485]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[329] ),
        .I4(\out[1431]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [849]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[849]_i_2 
       (.I0(\f_permutation_l_/round_in [1099]),
        .I1(\f_permutation_l_/round_in [1354]),
        .I2(\out[1590]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1483]),
        .I4(\out[1548]_i_16_n_0 ),
        .O(\out[849]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96699999)) 
    \out[84]_i_1 
       (.I0(\out[1262]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[619] ),
        .I2(\f_permutation_l_/out_reg_n_0_[210] ),
        .I3(\out[1598]_i_3_n_0 ),
        .I4(\out[276]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [84]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[850]_i_1 
       (.I0(\out[850]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[761] ),
        .I2(\out[1486]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[330] ),
        .I4(\out[1432]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [850]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[850]_i_2 
       (.I0(\f_permutation_l_/round_in [1100]),
        .I1(\f_permutation_l_/round_in [1355]),
        .I2(\out[1591]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1484]),
        .I4(\out[1549]_i_16_n_0 ),
        .O(\out[850]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[851]_i_1 
       (.I0(\out[851]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[762] ),
        .I2(\out[1487]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[331] ),
        .I4(\out[1433]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [851]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[851]_i_2 
       (.I0(\f_permutation_l_/round_in [1101]),
        .I1(\f_permutation_l_/round_in [1356]),
        .I2(\out[1592]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1485]),
        .I4(\out[1550]_i_16_n_0 ),
        .O(\out[851]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[852]_i_1 
       (.I0(\out[852]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[763] ),
        .I2(\out[1488]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[332] ),
        .I4(\out[1434]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [852]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[852]_i_2 
       (.I0(\f_permutation_l_/round_in [1102]),
        .I1(\f_permutation_l_/round_in [1357]),
        .I2(\out[1593]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1486]),
        .I4(\out[1551]_i_17_n_0 ),
        .O(\out[852]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[853]_i_1 
       (.I0(\out[853]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[764] ),
        .I2(\out[1489]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[333] ),
        .I4(\out[1435]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [853]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[853]_i_2 
       (.I0(\f_permutation_l_/round_in [1103]),
        .I1(\f_permutation_l_/round_in [1358]),
        .I2(\out[1594]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1487]),
        .I4(\out[1552]_i_16_n_0 ),
        .O(\out[853]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[854]_i_1 
       (.I0(\out[854]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[765] ),
        .I2(\out[1490]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[334] ),
        .I4(\out[1436]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [854]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[854]_i_2 
       (.I0(\f_permutation_l_/round_in [1104]),
        .I1(\f_permutation_l_/round_in [1359]),
        .I2(\out[1595]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1488]),
        .I4(\out[1553]_i_16_n_0 ),
        .O(\out[854]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[855]_i_1 
       (.I0(\out[855]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[766] ),
        .I2(\out[1491]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[335] ),
        .I4(\out[1437]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [855]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[855]_i_2 
       (.I0(\f_permutation_l_/round_in [1105]),
        .I1(\f_permutation_l_/round_in [1360]),
        .I2(\out[1596]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1489]),
        .I4(\out[1554]_i_16_n_0 ),
        .O(\out[855]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[856]_i_1 
       (.I0(\out[856]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[767] ),
        .I2(\out[1492]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[336] ),
        .I4(\out[1438]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [856]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[856]_i_2 
       (.I0(\f_permutation_l_/round_in [1106]),
        .I1(\f_permutation_l_/round_in [1361]),
        .I2(\out[1597]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1490]),
        .I4(\out[1555]_i_16_n_0 ),
        .O(\out[856]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[857]_i_1 
       (.I0(\out[857]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[704] ),
        .I2(\out[1493]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[337] ),
        .I4(\out[1439]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [857]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[857]_i_2 
       (.I0(\f_permutation_l_/round_in [1107]),
        .I1(\f_permutation_l_/round_in [1362]),
        .I2(\out[1598]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1491]),
        .I4(\out[1556]_i_16_n_0 ),
        .O(\out[857]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[858]_i_1 
       (.I0(\out[858]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[705] ),
        .I2(\out[1494]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[338] ),
        .I4(\out[1440]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [858]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[858]_i_2 
       (.I0(\f_permutation_l_/round_in [1108]),
        .I1(\f_permutation_l_/round_in [1363]),
        .I2(\out[1599]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1492]),
        .I4(\out[1557]_i_15_n_0 ),
        .O(\out[858]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[859]_i_1 
       (.I0(\out[859]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[706] ),
        .I2(\out[1495]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[339] ),
        .I4(\out[1441]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [859]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[859]_i_2 
       (.I0(\f_permutation_l_/round_in [1109]),
        .I1(\f_permutation_l_/round_in [1364]),
        .I2(\out[1536]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1493]),
        .I4(\out[1536]_i_14_n_0 ),
        .O(\out[859]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[85]_i_1 
       (.I0(\out[1263]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[620] ),
        .I2(\f_permutation_l_/out_reg_n_0_[211] ),
        .I3(\out[1343]_i_3_n_0 ),
        .I4(\out[277]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [85]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96AAAA96)) 
    \out[860]_i_1 
       (.I0(\out[860]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[707] ),
        .I2(\out[1496]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[340] ),
        .I4(\out[1442]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [860]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[860]_i_2 
       (.I0(\f_permutation_l_/round_in [1110]),
        .I1(\f_permutation_l_/round_in [1365]),
        .I2(\out[1537]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1494]),
        .I4(\out[1537]_i_10_n_0 ),
        .O(\out[860]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[861]_i_1 
       (.I0(\out[861]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[708] ),
        .I2(\out[1497]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[341] ),
        .I4(\out[1443]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [861]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[861]_i_2 
       (.I0(\f_permutation_l_/round_in [1111]),
        .I1(\f_permutation_l_/round_in [1366]),
        .I2(\out[1538]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1495]),
        .I4(\out[1538]_i_9_n_0 ),
        .O(\out[861]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[862]_i_1 
       (.I0(\out[926]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[709] ),
        .I2(\out[1498]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[342] ),
        .I4(\out[1444]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [862]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[863]_i_1 
       (.I0(\out[863]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[710] ),
        .I2(\out[1499]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[343] ),
        .I4(\out[1445]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [863]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[863]_i_2 
       (.I0(\f_permutation_l_/round_in [1113]),
        .I1(\f_permutation_l_/round_in [1368]),
        .I2(\out[1540]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1497]),
        .I4(\out[1540]_i_9_n_0 ),
        .O(\out[863]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[864]_i_1 
       (.I0(\out[864]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[711] ),
        .I2(\out[1500]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[344] ),
        .I4(\out[1446]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [864]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[864]_i_2 
       (.I0(\f_permutation_l_/round_in [1114]),
        .I1(\f_permutation_l_/round_in [1369]),
        .I2(\out[1541]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1498]),
        .I4(\out[1541]_i_9_n_0 ),
        .O(\out[864]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[865]_i_1 
       (.I0(\out[865]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[712] ),
        .I2(\out[1501]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[345] ),
        .I4(\out[1447]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [865]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[865]_i_2 
       (.I0(\f_permutation_l_/round_in [1115]),
        .I1(\f_permutation_l_/round_in [1370]),
        .I2(\out[1542]_i_12_n_0 ),
        .I3(\f_permutation_l_/round_in [1499]),
        .I4(\out[1542]_i_11_n_0 ),
        .O(\out[865]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[866]_i_1 
       (.I0(\out[866]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[713] ),
        .I2(\out[1502]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[346] ),
        .I4(\out[1448]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [866]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[866]_i_2 
       (.I0(\f_permutation_l_/round_in [1116]),
        .I1(\f_permutation_l_/round_in [1371]),
        .I2(\out[1543]_i_13_n_0 ),
        .I3(\f_permutation_l_/round_in [1500]),
        .I4(\out[1543]_i_11_n_0 ),
        .O(\out[866]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[867]_i_1 
       (.I0(\out[867]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[714] ),
        .I2(\out[1503]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[347] ),
        .I4(\out[1449]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [867]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[867]_i_2 
       (.I0(\f_permutation_l_/round_in [1117]),
        .I1(\f_permutation_l_/round_in [1372]),
        .I2(\out[1544]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1501]),
        .I4(\out[1544]_i_9_n_0 ),
        .O(\out[867]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[868]_i_1 
       (.I0(\out[868]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[715] ),
        .I2(\out[1504]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[348] ),
        .I4(\out[1450]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [868]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[868]_i_2 
       (.I0(\f_permutation_l_/round_in [1118]),
        .I1(\f_permutation_l_/round_in [1373]),
        .I2(\out[1545]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1502]),
        .I4(\out[1545]_i_9_n_0 ),
        .O(\out[868]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[869]_i_1 
       (.I0(\out[869]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[716] ),
        .I2(\out[1505]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[349] ),
        .I4(\out[1451]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [869]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[869]_i_2 
       (.I0(\f_permutation_l_/round_in [1119]),
        .I1(\f_permutation_l_/round_in [1374]),
        .I2(\out[1546]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1503]),
        .I4(\out[1546]_i_9_n_0 ),
        .O(\out[869]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[86]_i_1 
       (.I0(\out[1264]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[621] ),
        .I2(\f_permutation_l_/out_reg_n_0_[212] ),
        .I3(\out[1280]_i_3_n_0 ),
        .I4(\out[278]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [86]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[870]_i_1 
       (.I0(\out[870]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[717] ),
        .I2(\out[1506]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[350] ),
        .I4(\out[1452]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [870]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[870]_i_2 
       (.I0(\f_permutation_l_/round_in [1120]),
        .I1(\f_permutation_l_/round_in [1375]),
        .I2(\out[1547]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1504]),
        .I4(\out[1547]_i_9_n_0 ),
        .O(\out[870]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[871]_i_1 
       (.I0(\out[871]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[718] ),
        .I2(\out[1507]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[351] ),
        .I4(\out[1453]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [871]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[871]_i_2 
       (.I0(\f_permutation_l_/round_in [1121]),
        .I1(\f_permutation_l_/round_in [1376]),
        .I2(\out[1548]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1505]),
        .I4(\out[1548]_i_9_n_0 ),
        .O(\out[871]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[872]_i_1 
       (.I0(\out[872]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[719] ),
        .I2(\out[1508]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[352] ),
        .I4(\out[1454]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [872]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[872]_i_2 
       (.I0(\f_permutation_l_/round_in [1122]),
        .I1(\f_permutation_l_/round_in [1377]),
        .I2(\out[1549]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1506]),
        .I4(\out[1549]_i_9_n_0 ),
        .O(\out[872]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[873]_i_1 
       (.I0(\out[873]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[720] ),
        .I2(\out[1509]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[353] ),
        .I4(\out[1455]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [873]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[873]_i_2 
       (.I0(\f_permutation_l_/round_in [1123]),
        .I1(\f_permutation_l_/round_in [1378]),
        .I2(\out[1550]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1507]),
        .I4(\out[1550]_i_9_n_0 ),
        .O(\out[873]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[874]_i_1 
       (.I0(\out[874]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[721] ),
        .I2(\out[1510]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[354] ),
        .I4(\out[1456]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [874]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[874]_i_2 
       (.I0(\f_permutation_l_/round_in [1124]),
        .I1(\f_permutation_l_/round_in [1379]),
        .I2(\out[1551]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1508]),
        .I4(\out[1551]_i_10_n_0 ),
        .O(\out[874]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[875]_i_1 
       (.I0(\out[875]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[722] ),
        .I2(\out[1511]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[355] ),
        .I4(\out[1457]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [875]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[875]_i_2 
       (.I0(\f_permutation_l_/round_in [1125]),
        .I1(\f_permutation_l_/round_in [1380]),
        .I2(\out[1552]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1509]),
        .I4(\out[1552]_i_9_n_0 ),
        .O(\out[875]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[876]_i_1 
       (.I0(\out[876]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[723] ),
        .I2(\out[1512]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[356] ),
        .I4(\out[1458]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [876]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[876]_i_2 
       (.I0(\f_permutation_l_/round_in [1126]),
        .I1(\f_permutation_l_/round_in [1381]),
        .I2(\out[1553]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1510]),
        .I4(\out[1553]_i_9_n_0 ),
        .O(\out[876]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[877]_i_1 
       (.I0(\out[877]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[724] ),
        .I2(\out[1513]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[357] ),
        .I4(\out[1459]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [877]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[877]_i_2 
       (.I0(\f_permutation_l_/round_in [1127]),
        .I1(\f_permutation_l_/round_in [1382]),
        .I2(\out[1554]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1511]),
        .I4(\out[1554]_i_9_n_0 ),
        .O(\out[877]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[878]_i_1 
       (.I0(\out[878]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[725] ),
        .I2(\out[1514]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[358] ),
        .I4(\out[1460]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [878]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[878]_i_2 
       (.I0(\f_permutation_l_/round_in [1128]),
        .I1(\f_permutation_l_/round_in [1383]),
        .I2(\out[1555]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1512]),
        .I4(\out[1555]_i_9_n_0 ),
        .O(\out[878]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA6969AA)) 
    \out[879]_i_1 
       (.I0(\out[879]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[726] ),
        .I2(\out[1515]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[359] ),
        .I4(\out[1461]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [879]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[879]_i_2 
       (.I0(\f_permutation_l_/round_in [1129]),
        .I1(\f_permutation_l_/round_in [1384]),
        .I2(\out[1556]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1513]),
        .I4(\out[1556]_i_10_n_0 ),
        .O(\out[879]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[87]_i_1 
       (.I0(\out[1265]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[622] ),
        .I2(\f_permutation_l_/out_reg_n_0_[213] ),
        .I3(\out[1281]_i_3_n_0 ),
        .I4(\out[279]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [87]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[880]_i_1 
       (.I0(\out[880]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[727] ),
        .I2(\out[1516]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[360] ),
        .I4(\out[1462]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [880]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[880]_i_2 
       (.I0(\f_permutation_l_/round_in [1130]),
        .I1(\f_permutation_l_/round_in [1385]),
        .I2(\out[1557]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1514]),
        .I4(\out[1557]_i_9_n_0 ),
        .O(\out[880]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[881]_i_1 
       (.I0(\out[881]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[728] ),
        .I2(\out[1517]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[361] ),
        .I4(\out[1463]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [881]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[881]_i_2 
       (.I0(\f_permutation_l_/round_in [1131]),
        .I1(\f_permutation_l_/round_in [1386]),
        .I2(\out[1558]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1515]),
        .I4(\out[1558]_i_9_n_0 ),
        .O(\out[881]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[882]_i_1 
       (.I0(\out[882]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[729] ),
        .I2(\out[1518]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[362] ),
        .I4(\out[1464]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [882]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[882]_i_2 
       (.I0(\f_permutation_l_/round_in [1132]),
        .I1(\f_permutation_l_/round_in [1387]),
        .I2(\out[1559]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1516]),
        .I4(\out[1559]_i_9_n_0 ),
        .O(\out[882]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[883]_i_1 
       (.I0(\out[883]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[730] ),
        .I2(\out[1519]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[363] ),
        .I4(\out[1465]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [883]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[883]_i_2 
       (.I0(\f_permutation_l_/round_in [1133]),
        .I1(\f_permutation_l_/round_in [1388]),
        .I2(\out[1560]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1517]),
        .I4(\out[1560]_i_9_n_0 ),
        .O(\out[883]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[884]_i_1 
       (.I0(\out[884]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[731] ),
        .I2(\out[1520]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[364] ),
        .I4(\out[1466]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [884]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[884]_i_2 
       (.I0(\f_permutation_l_/round_in [1134]),
        .I1(\f_permutation_l_/round_in [1389]),
        .I2(\out[1561]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1518]),
        .I4(\out[1561]_i_9_n_0 ),
        .O(\out[884]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[885]_i_1 
       (.I0(\out[885]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[732] ),
        .I2(\out[1521]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[365] ),
        .I4(\out[1467]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [885]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[885]_i_2 
       (.I0(\f_permutation_l_/round_in [1135]),
        .I1(\f_permutation_l_/round_in [1390]),
        .I2(\out[1562]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1519]),
        .I4(\out[1562]_i_9_n_0 ),
        .O(\out[885]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[886]_i_1 
       (.I0(\out[886]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[733] ),
        .I2(\out[1522]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[366] ),
        .I4(\out[1468]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [886]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[886]_i_2 
       (.I0(\f_permutation_l_/round_in [1136]),
        .I1(\f_permutation_l_/round_in [1391]),
        .I2(\out[1563]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1520]),
        .I4(\out[1563]_i_9_n_0 ),
        .O(\out[886]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[887]_i_1 
       (.I0(\out[887]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[734] ),
        .I2(\out[1523]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[367] ),
        .I4(\out[1469]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [887]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[887]_i_2 
       (.I0(\f_permutation_l_/round_in [1137]),
        .I1(\f_permutation_l_/round_in [1392]),
        .I2(\out[1564]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1521]),
        .I4(\out[1564]_i_9_n_0 ),
        .O(\out[887]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[888]_i_1 
       (.I0(\out[888]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[735] ),
        .I2(\out[1524]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[368] ),
        .I4(\out[1470]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [888]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[888]_i_2 
       (.I0(\f_permutation_l_/round_in [1138]),
        .I1(\f_permutation_l_/round_in [1393]),
        .I2(\out[1565]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1522]),
        .I4(\out[1565]_i_9_n_0 ),
        .O(\out[888]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[889]_i_1 
       (.I0(\out[889]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[736] ),
        .I2(\out[1525]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[369] ),
        .I4(\out[1471]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [889]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[889]_i_2 
       (.I0(\f_permutation_l_/round_in [1139]),
        .I1(\f_permutation_l_/round_in [1394]),
        .I2(\out[1566]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1523]),
        .I4(\out[1566]_i_9_n_0 ),
        .O(\out[889]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[88]_i_1 
       (.I0(\out[1266]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[623] ),
        .I2(\f_permutation_l_/out_reg_n_0_[214] ),
        .I3(\out[1538]_i_3_n_0 ),
        .I4(\out[280]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [88]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[890]_i_1 
       (.I0(\out[890]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[737] ),
        .I2(\out[1526]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[370] ),
        .I4(\out[1408]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [890]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[890]_i_2 
       (.I0(\f_permutation_l_/round_in [1140]),
        .I1(\f_permutation_l_/round_in [1395]),
        .I2(\out[1567]_i_11_n_0 ),
        .I3(\f_permutation_l_/round_in [1524]),
        .I4(\out[1567]_i_10_n_0 ),
        .O(\out[890]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[891]_i_1 
       (.I0(\out[891]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[738] ),
        .I2(\out[1527]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[371] ),
        .I4(\out[1409]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [891]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[891]_i_2 
       (.I0(\f_permutation_l_/round_in [1141]),
        .I1(\f_permutation_l_/round_in [1396]),
        .I2(\out[1568]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1525]),
        .I4(\out[1568]_i_9_n_0 ),
        .O(\out[891]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[892]_i_1 
       (.I0(\out[892]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[739] ),
        .I2(\out[1528]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[372] ),
        .I4(\out[1410]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [892]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[892]_i_2 
       (.I0(\f_permutation_l_/round_in [1142]),
        .I1(\f_permutation_l_/round_in [1397]),
        .I2(\out[1569]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1526]),
        .I4(\out[1569]_i_9_n_0 ),
        .O(\out[892]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[893]_i_1 
       (.I0(\out[893]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[740] ),
        .I2(\out[1529]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[373] ),
        .I4(\out[1411]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [893]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[893]_i_2 
       (.I0(\f_permutation_l_/round_in [1143]),
        .I1(\f_permutation_l_/round_in [1398]),
        .I2(\out[1570]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1527]),
        .I4(\out[1570]_i_9_n_0 ),
        .O(\out[893]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[894]_i_1 
       (.I0(\out[894]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[741] ),
        .I2(\out[1530]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[374] ),
        .I4(\out[1412]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [894]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[894]_i_2 
       (.I0(\f_permutation_l_/round_in [1144]),
        .I1(\f_permutation_l_/round_in [1399]),
        .I2(\out[1571]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1528]),
        .I4(\out[1571]_i_9_n_0 ),
        .O(\out[894]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAA9696AA)) 
    \out[895]_i_1 
       (.I0(\out[895]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[742] ),
        .I2(\out[1531]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[375] ),
        .I4(\out[1413]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [895]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[895]_i_2 
       (.I0(\f_permutation_l_/round_in [1145]),
        .I1(\f_permutation_l_/round_in [1400]),
        .I2(\out[1572]_i_10_n_0 ),
        .I3(\f_permutation_l_/round_in [1529]),
        .I4(\out[1572]_i_9_n_0 ),
        .O(\out[895]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[896]_i_1 
       (.I0(\f_permutation_l_/round_in [1146]),
        .I1(\out[1573]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[743] ),
        .I3(\out[1532]_i_3_n_0 ),
        .I4(\out[896]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [896]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[896]_i_2 
       (.I0(padder_out_1[66]),
        .I1(out[2]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1146]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[896]_i_3 
       (.I0(\f_permutation_l_/round_in [1535]),
        .I1(\f_permutation_l_/round_in [1470]),
        .I2(\out[1579]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1599]),
        .I4(\out[1579]_i_7_n_0 ),
        .O(\out[896]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[897]_i_1 
       (.I0(\f_permutation_l_/round_in [1147]),
        .I1(\out[1574]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[744] ),
        .I3(\out[1533]_i_3_n_0 ),
        .I4(\out[897]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [897]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[897]_i_2 
       (.I0(padder_out_1[67]),
        .I1(out[3]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1147]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[897]_i_3 
       (.I0(\f_permutation_l_/round_in [1472]),
        .I1(\f_permutation_l_/round_in [1471]),
        .I2(\out[1580]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1536]),
        .I4(\out[1580]_i_6_n_0 ),
        .O(\out[897]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[898]_i_1 
       (.I0(\f_permutation_l_/round_in [1148]),
        .I1(\out[1575]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[745] ),
        .I3(\out[1534]_i_3_n_0 ),
        .I4(\out[898]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [898]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[898]_i_2 
       (.I0(padder_out_1[68]),
        .I1(out[4]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1148]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[898]_i_3 
       (.I0(\f_permutation_l_/round_in [1473]),
        .I1(\f_permutation_l_/round_in [1408]),
        .I2(\out[1581]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1537]),
        .I4(\out[1581]_i_6_n_0 ),
        .O(\out[898]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[899]_i_1 
       (.I0(\f_permutation_l_/round_in [1149]),
        .I1(\out[1576]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[746] ),
        .I3(\out[1535]_i_2_n_0 ),
        .I4(\out[899]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [899]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[899]_i_2 
       (.I0(padder_out_1[69]),
        .I1(out[5]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1149]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[899]_i_3 
       (.I0(\f_permutation_l_/round_in [1474]),
        .I1(\f_permutation_l_/round_in [1409]),
        .I2(\out[1582]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1538]),
        .I4(\out[1582]_i_6_n_0 ),
        .O(\out[899]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[89]_i_1 
       (.I0(\out[1267]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[624] ),
        .I2(\f_permutation_l_/out_reg_n_0_[215] ),
        .I3(\out[1539]_i_3_n_0 ),
        .I4(\out[281]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [89]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96999996)) 
    \out[8]_i_1 
       (.I0(\out[1586]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[198] ),
        .I2(\out[264]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1041]),
        .I4(\out[1510]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[900]_i_1 
       (.I0(\f_permutation_l_/round_in [1150]),
        .I1(\out[1577]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[747] ),
        .I3(\out[1472]_i_3_n_0 ),
        .I4(\out[900]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [900]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[900]_i_2 
       (.I0(padder_out_1[70]),
        .I1(out[6]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1150]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[900]_i_3 
       (.I0(\f_permutation_l_/round_in [1475]),
        .I1(\f_permutation_l_/round_in [1410]),
        .I2(\out[1583]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1539]),
        .I4(\out[1583]_i_6_n_0 ),
        .O(\out[900]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[901]_i_1 
       (.I0(\f_permutation_l_/round_in [1151]),
        .I1(\out[1578]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[748] ),
        .I3(\out[1473]_i_2_n_0 ),
        .I4(\out[901]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [901]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[901]_i_2 
       (.I0(padder_out_1[71]),
        .I1(out[7]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1151]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[901]_i_3 
       (.I0(\f_permutation_l_/round_in [1476]),
        .I1(\f_permutation_l_/round_in [1411]),
        .I2(\out[1584]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1540]),
        .I4(\out[1584]_i_6_n_0 ),
        .O(\out[901]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[902]_i_1 
       (.I0(\f_permutation_l_/round_in [1088]),
        .I1(\out[1579]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[749] ),
        .I3(\out[1474]_i_3_n_0 ),
        .I4(\out[902]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [902]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[902]_i_2 
       (.I0(padder_out_1[120]),
        .I1(out[56]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1088]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[902]_i_3 
       (.I0(\f_permutation_l_/round_in [1477]),
        .I1(\f_permutation_l_/round_in [1412]),
        .I2(\out[1585]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1541]),
        .I4(\out[1585]_i_6_n_0 ),
        .O(\out[902]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[903]_i_1 
       (.I0(\f_permutation_l_/round_in [1089]),
        .I1(\out[1580]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[750] ),
        .I3(\out[1475]_i_2_n_0 ),
        .I4(\out[903]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [903]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[903]_i_2 
       (.I0(padder_out_1[121]),
        .I1(out[57]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1089]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[903]_i_3 
       (.I0(\f_permutation_l_/round_in [1478]),
        .I1(\f_permutation_l_/round_in [1413]),
        .I2(\out[1586]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1542]),
        .I4(\out[1586]_i_6_n_0 ),
        .O(\out[903]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[904]_i_1 
       (.I0(\f_permutation_l_/round_in [1090]),
        .I1(\out[1581]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[751] ),
        .I3(\out[1476]_i_3_n_0 ),
        .I4(\out[904]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [904]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[904]_i_2 
       (.I0(padder_out_1[122]),
        .I1(out[58]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1090]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[904]_i_3 
       (.I0(\f_permutation_l_/round_in [1479]),
        .I1(\f_permutation_l_/round_in [1414]),
        .I2(\out[1587]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1543]),
        .I4(\out[1587]_i_6_n_0 ),
        .O(\out[904]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[905]_i_1 
       (.I0(\f_permutation_l_/round_in [1091]),
        .I1(\out[1582]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[752] ),
        .I3(\out[1477]_i_3_n_0 ),
        .I4(\out[905]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [905]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[905]_i_2 
       (.I0(padder_out_1[123]),
        .I1(out[59]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1091]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[905]_i_3 
       (.I0(\f_permutation_l_/round_in [1480]),
        .I1(\f_permutation_l_/round_in [1415]),
        .I2(\out[1588]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1544]),
        .I4(\out[1588]_i_6_n_0 ),
        .O(\out[905]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[906]_i_1 
       (.I0(\f_permutation_l_/round_in [1092]),
        .I1(\out[1583]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[753] ),
        .I3(\out[1478]_i_3_n_0 ),
        .I4(\out[906]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [906]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[906]_i_2 
       (.I0(padder_out_1[124]),
        .I1(out[60]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1092]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[906]_i_3 
       (.I0(\f_permutation_l_/round_in [1481]),
        .I1(\f_permutation_l_/round_in [1416]),
        .I2(\out[1589]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1545]),
        .I4(\out[1589]_i_6_n_0 ),
        .O(\out[906]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[907]_i_1 
       (.I0(\f_permutation_l_/round_in [1093]),
        .I1(\out[1584]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[754] ),
        .I3(\out[1479]_i_2_n_0 ),
        .I4(\out[907]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [907]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[907]_i_2 
       (.I0(padder_out_1[125]),
        .I1(out[61]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1093]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[907]_i_3 
       (.I0(\f_permutation_l_/round_in [1482]),
        .I1(\f_permutation_l_/round_in [1417]),
        .I2(\out[1590]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1546]),
        .I4(\out[1590]_i_6_n_0 ),
        .O(\out[907]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[908]_i_1 
       (.I0(\f_permutation_l_/round_in [1094]),
        .I1(\out[1585]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[755] ),
        .I3(\out[1480]_i_3_n_0 ),
        .I4(\out[908]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [908]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[908]_i_2 
       (.I0(padder_out_1[126]),
        .I1(out[62]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1094]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[908]_i_3 
       (.I0(\f_permutation_l_/round_in [1483]),
        .I1(\f_permutation_l_/round_in [1418]),
        .I2(\out[1591]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1547]),
        .I4(\out[1591]_i_6_n_0 ),
        .O(\out[908]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[909]_i_1 
       (.I0(\f_permutation_l_/round_in [1095]),
        .I1(\out[1586]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[756] ),
        .I3(\out[1481]_i_3_n_0 ),
        .I4(\out[909]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [909]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[909]_i_2 
       (.I0(padder_out_1[127]),
        .I1(out[63]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1095]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[909]_i_3 
       (.I0(\f_permutation_l_/round_in [1484]),
        .I1(\f_permutation_l_/round_in [1419]),
        .I2(\out[1592]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1548]),
        .I4(\out[1592]_i_6_n_0 ),
        .O(\out[909]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[90]_i_1 
       (.I0(\out[1268]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[625] ),
        .I2(\f_permutation_l_/out_reg_n_0_[216] ),
        .I3(\out[1540]_i_3_n_0 ),
        .I4(\out[282]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [90]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[910]_i_1 
       (.I0(\f_permutation_l_/round_in [1096]),
        .I1(\out[1587]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[757] ),
        .I3(\out[1482]_i_3_n_0 ),
        .I4(\out[910]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [910]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[910]_i_2 
       (.I0(padder_out_1[112]),
        .I1(out[48]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1096]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[910]_i_3 
       (.I0(\f_permutation_l_/round_in [1485]),
        .I1(\f_permutation_l_/round_in [1420]),
        .I2(\out[1593]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1549]),
        .I4(\out[1593]_i_6_n_0 ),
        .O(\out[910]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[911]_i_1 
       (.I0(\f_permutation_l_/round_in [1097]),
        .I1(\out[1588]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[758] ),
        .I3(\out[1483]_i_3_n_0 ),
        .I4(\out[911]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [911]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[911]_i_2 
       (.I0(padder_out_1[113]),
        .I1(out[49]),
        .I2(\out[911]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1097]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[911]_i_3 
       (.I0(\f_permutation_l_/round_in [1486]),
        .I1(\f_permutation_l_/round_in [1421]),
        .I2(\out[1594]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1550]),
        .I4(\out[1594]_i_6_n_0 ),
        .O(\out[911]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \out[911]_i_4 
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(\out[911]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[912]_i_1 
       (.I0(\f_permutation_l_/round_in [1098]),
        .I1(\out[1589]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[759] ),
        .I3(\out[1484]_i_3_n_0 ),
        .I4(\out[912]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [912]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[912]_i_2 
       (.I0(padder_out_1[114]),
        .I1(out[50]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1098]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[912]_i_3 
       (.I0(\f_permutation_l_/round_in [1487]),
        .I1(\f_permutation_l_/round_in [1422]),
        .I2(\out[1595]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1551]),
        .I4(\out[1595]_i_6_n_0 ),
        .O(\out[912]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[913]_i_1 
       (.I0(\f_permutation_l_/round_in [1099]),
        .I1(\out[1590]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[760] ),
        .I3(\out[1485]_i_3_n_0 ),
        .I4(\out[913]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [913]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[913]_i_2 
       (.I0(padder_out_1[115]),
        .I1(out[51]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1099]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[913]_i_3 
       (.I0(\f_permutation_l_/round_in [1488]),
        .I1(\f_permutation_l_/round_in [1423]),
        .I2(\out[1596]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1552]),
        .I4(\out[1596]_i_6_n_0 ),
        .O(\out[913]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[914]_i_1 
       (.I0(\f_permutation_l_/round_in [1100]),
        .I1(\out[1591]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[761] ),
        .I3(\out[1486]_i_3_n_0 ),
        .I4(\out[914]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [914]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[914]_i_2 
       (.I0(padder_out_1[116]),
        .I1(out[52]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1100]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[914]_i_3 
       (.I0(\f_permutation_l_/round_in [1489]),
        .I1(\f_permutation_l_/round_in [1424]),
        .I2(\out[1597]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1553]),
        .I4(\out[1597]_i_6_n_0 ),
        .O(\out[914]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[915]_i_1 
       (.I0(\f_permutation_l_/round_in [1101]),
        .I1(\out[1592]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[762] ),
        .I3(\out[1487]_i_2_n_0 ),
        .I4(\out[915]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [915]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[915]_i_2 
       (.I0(padder_out_1[117]),
        .I1(out[53]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1101]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[915]_i_3 
       (.I0(\f_permutation_l_/round_in [1490]),
        .I1(\f_permutation_l_/round_in [1425]),
        .I2(\out[1598]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1554]),
        .I4(\out[1598]_i_6_n_0 ),
        .O(\out[915]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[916]_i_1 
       (.I0(\f_permutation_l_/round_in [1102]),
        .I1(\out[1593]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[763] ),
        .I3(\out[1488]_i_3_n_0 ),
        .I4(\out[916]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [916]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[916]_i_2 
       (.I0(padder_out_1[118]),
        .I1(out[54]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1102]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[916]_i_3 
       (.I0(\f_permutation_l_/round_in [1491]),
        .I1(\f_permutation_l_/round_in [1426]),
        .I2(\out[1599]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1555]),
        .I4(\out[1599]_i_8_n_0 ),
        .O(\out[916]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[917]_i_1 
       (.I0(\f_permutation_l_/round_in [1103]),
        .I1(\out[1594]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[764] ),
        .I3(\out[1489]_i_3_n_0 ),
        .I4(\out[917]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [917]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[917]_i_2 
       (.I0(padder_out_1[119]),
        .I1(out[55]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1103]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[917]_i_3 
       (.I0(\f_permutation_l_/round_in [1492]),
        .I1(\f_permutation_l_/round_in [1427]),
        .I2(\out[1536]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1556]),
        .I4(\out[1536]_i_10_n_0 ),
        .O(\out[917]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[918]_i_1 
       (.I0(\f_permutation_l_/round_in [1104]),
        .I1(\out[1595]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[765] ),
        .I3(\out[1490]_i_3_n_0 ),
        .I4(\out[918]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [918]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[918]_i_2 
       (.I0(padder_out_1[104]),
        .I1(out[40]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1104]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[918]_i_3 
       (.I0(\f_permutation_l_/round_in [1493]),
        .I1(\f_permutation_l_/round_in [1428]),
        .I2(\out[1537]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1557]),
        .I4(\out[1537]_i_9_n_0 ),
        .O(\out[918]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[919]_i_1 
       (.I0(\f_permutation_l_/round_in [1105]),
        .I1(\out[1596]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[766] ),
        .I3(\out[1491]_i_3_n_0 ),
        .I4(\out[919]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [919]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[919]_i_2 
       (.I0(padder_out_1[105]),
        .I1(out[41]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1105]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[919]_i_3 
       (.I0(\f_permutation_l_/round_in [1494]),
        .I1(\f_permutation_l_/round_in [1429]),
        .I2(\out[1538]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1558]),
        .I4(\out[1538]_i_6_n_0 ),
        .O(\out[919]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[91]_i_1 
       (.I0(\out[1269]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[626] ),
        .I2(\f_permutation_l_/out_reg_n_0_[217] ),
        .I3(\out[1541]_i_3_n_0 ),
        .I4(\out[283]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [91]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[920]_i_1 
       (.I0(\f_permutation_l_/round_in [1106]),
        .I1(\out[1597]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[767] ),
        .I3(\out[1492]_i_3_n_0 ),
        .I4(\out[920]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [920]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[920]_i_2 
       (.I0(padder_out_1[106]),
        .I1(out[42]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1106]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[920]_i_3 
       (.I0(\f_permutation_l_/round_in [1495]),
        .I1(\f_permutation_l_/round_in [1430]),
        .I2(\out[1539]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1559]),
        .I4(\out[1539]_i_8_n_0 ),
        .O(\out[920]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[921]_i_1 
       (.I0(\f_permutation_l_/round_in [1107]),
        .I1(\out[1598]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[704] ),
        .I3(\out[1493]_i_3_n_0 ),
        .I4(\out[921]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [921]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[921]_i_2 
       (.I0(padder_out_1[107]),
        .I1(out[43]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1107]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[921]_i_3 
       (.I0(\f_permutation_l_/round_in [1496]),
        .I1(\f_permutation_l_/round_in [1431]),
        .I2(\out[1540]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1560]),
        .I4(\out[1540]_i_6_n_0 ),
        .O(\out[921]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[922]_i_1 
       (.I0(\f_permutation_l_/round_in [1108]),
        .I1(\out[1599]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[705] ),
        .I3(\out[1494]_i_3_n_0 ),
        .I4(\out[922]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [922]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[922]_i_2 
       (.I0(padder_out_1[108]),
        .I1(out[44]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1108]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[922]_i_3 
       (.I0(\f_permutation_l_/round_in [1497]),
        .I1(\f_permutation_l_/round_in [1432]),
        .I2(\out[1541]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1561]),
        .I4(\out[1541]_i_6_n_0 ),
        .O(\out[922]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h6FF69009)) 
    \out[923]_i_1 
       (.I0(\f_permutation_l_/round_in [1109]),
        .I1(\out[1472]_i_2_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[706] ),
        .I3(\out[1495]_i_3_n_0 ),
        .I4(\out[923]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [923]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[923]_i_2 
       (.I0(padder_out_1[109]),
        .I1(out[45]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1109]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[923]_i_3 
       (.I0(\f_permutation_l_/round_in [1498]),
        .I1(\f_permutation_l_/round_in [1433]),
        .I2(\out[1542]_i_9_n_0 ),
        .I3(\f_permutation_l_/round_in [1562]),
        .I4(\out[1542]_i_7_n_0 ),
        .O(\out[923]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[924]_i_1 
       (.I0(\f_permutation_l_/round_in [1110]),
        .I1(\out[1537]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[707] ),
        .I3(\out[1496]_i_3_n_0 ),
        .I4(\out[924]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [924]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[924]_i_2 
       (.I0(padder_out_1[110]),
        .I1(out[46]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1110]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[924]_i_3 
       (.I0(\f_permutation_l_/round_in [1499]),
        .I1(\f_permutation_l_/round_in [1434]),
        .I2(\out[1543]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1563]),
        .I4(\out[1543]_i_10_n_0 ),
        .O(\out[924]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[925]_i_1 
       (.I0(\f_permutation_l_/round_in [1111]),
        .I1(\out[1538]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[708] ),
        .I3(\out[1497]_i_3_n_0 ),
        .I4(\out[925]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [925]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[925]_i_2 
       (.I0(padder_out_1[111]),
        .I1(out[47]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1111]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[925]_i_3 
       (.I0(\f_permutation_l_/round_in [1500]),
        .I1(\f_permutation_l_/round_in [1435]),
        .I2(\out[1544]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1564]),
        .I4(\out[1544]_i_6_n_0 ),
        .O(\out[925]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h41BEBE41)) 
    \out[926]_i_1 
       (.I0(\out[926]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[709] ),
        .I2(\out[1498]_i_3_n_0 ),
        .I3(\out[1545]_i_3_n_0 ),
        .I4(\f_permutation_l_/round_in [1501]),
        .O(\f_permutation_l_/round_out [926]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[926]_i_2 
       (.I0(\f_permutation_l_/round_in [1112]),
        .I1(\out[1539]_i_12_n_0 ),
        .I2(\f_permutation_l_/round_in [1367]),
        .I3(\f_permutation_l_/round_in [1496]),
        .I4(\out[1539]_i_14_n_0 ),
        .O(\out[926]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[926]_i_3 
       (.I0(padder_out_1[485]),
        .I1(out[421]),
        .I2(\out[1447]_i_4_n_0 ),
        .O(\f_permutation_l_/round_in [1501]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[926]_i_4 
       (.I0(padder_out_1[96]),
        .I1(out[32]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1112]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[927]_i_1 
       (.I0(\f_permutation_l_/round_in [1113]),
        .I1(\out[1540]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[710] ),
        .I3(\out[1499]_i_3_n_0 ),
        .I4(\out[927]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [927]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[927]_i_2 
       (.I0(padder_out_1[97]),
        .I1(out[33]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1113]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[927]_i_3 
       (.I0(\f_permutation_l_/round_in [1502]),
        .I1(\f_permutation_l_/round_in [1437]),
        .I2(\out[1546]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1566]),
        .I4(\out[1546]_i_6_n_0 ),
        .O(\out[927]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[928]_i_1 
       (.I0(\f_permutation_l_/round_in [1114]),
        .I1(\out[1541]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[711] ),
        .I3(\out[1500]_i_3_n_0 ),
        .I4(\out[928]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [928]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[928]_i_2 
       (.I0(padder_out_1[98]),
        .I1(out[34]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1114]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[928]_i_3 
       (.I0(\f_permutation_l_/round_in [1503]),
        .I1(\f_permutation_l_/round_in [1438]),
        .I2(\out[1547]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1567]),
        .I4(\out[1547]_i_6_n_0 ),
        .O(\out[928]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[929]_i_1 
       (.I0(\f_permutation_l_/round_in [1115]),
        .I1(\out[1542]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[712] ),
        .I3(\out[1501]_i_3_n_0 ),
        .I4(\out[929]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [929]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[929]_i_2 
       (.I0(padder_out_1[99]),
        .I1(out[35]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1115]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[929]_i_3 
       (.I0(\f_permutation_l_/round_in [1504]),
        .I1(\f_permutation_l_/round_in [1439]),
        .I2(\out[1548]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1568]),
        .I4(\out[1548]_i_6_n_0 ),
        .O(\out[929]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[92]_i_1 
       (.I0(\out[1270]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[627] ),
        .I2(\f_permutation_l_/out_reg_n_0_[218] ),
        .I3(\out[1542]_i_3_n_0 ),
        .I4(\out[284]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [92]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[930]_i_1 
       (.I0(\f_permutation_l_/round_in [1116]),
        .I1(\out[1543]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[713] ),
        .I3(\out[1502]_i_3_n_0 ),
        .I4(\out[930]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [930]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[930]_i_2 
       (.I0(padder_out_1[100]),
        .I1(out[36]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1116]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[930]_i_3 
       (.I0(\f_permutation_l_/round_in [1505]),
        .I1(\f_permutation_l_/round_in [1440]),
        .I2(\out[1549]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1569]),
        .I4(\out[1549]_i_6_n_0 ),
        .O(\out[930]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[931]_i_1 
       (.I0(\f_permutation_l_/round_in [1117]),
        .I1(\out[1544]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[714] ),
        .I3(\out[1503]_i_2_n_0 ),
        .I4(\out[931]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [931]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[931]_i_2 
       (.I0(padder_out_1[101]),
        .I1(out[37]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1117]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[931]_i_3 
       (.I0(\f_permutation_l_/round_in [1506]),
        .I1(\f_permutation_l_/round_in [1441]),
        .I2(\out[1550]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1570]),
        .I4(\out[1550]_i_6_n_0 ),
        .O(\out[931]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[932]_i_1 
       (.I0(\f_permutation_l_/round_in [1118]),
        .I1(\out[1545]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[715] ),
        .I3(\out[1504]_i_3_n_0 ),
        .I4(\out[932]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [932]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[932]_i_2 
       (.I0(padder_out_1[102]),
        .I1(out[38]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1118]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[932]_i_3 
       (.I0(\f_permutation_l_/round_in [1507]),
        .I1(\f_permutation_l_/round_in [1442]),
        .I2(\out[1551]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1571]),
        .I4(\out[1551]_i_9_n_0 ),
        .O(\out[932]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[933]_i_1 
       (.I0(\f_permutation_l_/round_in [1119]),
        .I1(\out[1546]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[716] ),
        .I3(\out[1505]_i_3_n_0 ),
        .I4(\out[933]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [933]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[933]_i_2 
       (.I0(padder_out_1[103]),
        .I1(out[39]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1119]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[933]_i_3 
       (.I0(\f_permutation_l_/round_in [1508]),
        .I1(\f_permutation_l_/round_in [1443]),
        .I2(\out[1552]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1572]),
        .I4(\out[1552]_i_6_n_0 ),
        .O(\out[933]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[934]_i_1 
       (.I0(\f_permutation_l_/round_in [1120]),
        .I1(\out[1547]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[717] ),
        .I3(\out[1506]_i_3_n_0 ),
        .I4(\out[934]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [934]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[934]_i_2 
       (.I0(padder_out_1[88]),
        .I1(out[24]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1120]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[934]_i_3 
       (.I0(\f_permutation_l_/round_in [1509]),
        .I1(\f_permutation_l_/round_in [1444]),
        .I2(\out[1553]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1573]),
        .I4(\out[1553]_i_6_n_0 ),
        .O(\out[934]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[935]_i_1 
       (.I0(\f_permutation_l_/round_in [1121]),
        .I1(\out[1548]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[718] ),
        .I3(\out[1507]_i_3_n_0 ),
        .I4(\out[935]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [935]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[935]_i_2 
       (.I0(padder_out_1[89]),
        .I1(out[25]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1121]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[935]_i_3 
       (.I0(\f_permutation_l_/round_in [1510]),
        .I1(\f_permutation_l_/round_in [1445]),
        .I2(\out[1554]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1574]),
        .I4(\out[1554]_i_6_n_0 ),
        .O(\out[935]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[936]_i_1 
       (.I0(\f_permutation_l_/round_in [1122]),
        .I1(\out[1549]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[719] ),
        .I3(\out[1508]_i_3_n_0 ),
        .I4(\out[936]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [936]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[936]_i_2 
       (.I0(padder_out_1[90]),
        .I1(out[26]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1122]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[936]_i_3 
       (.I0(\f_permutation_l_/round_in [1511]),
        .I1(\f_permutation_l_/round_in [1446]),
        .I2(\out[1555]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1575]),
        .I4(\out[1555]_i_6_n_0 ),
        .O(\out[936]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[937]_i_1 
       (.I0(\f_permutation_l_/round_in [1123]),
        .I1(\out[1550]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[720] ),
        .I3(\out[1509]_i_3_n_0 ),
        .I4(\out[937]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [937]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[937]_i_2 
       (.I0(padder_out_1[91]),
        .I1(out[27]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1123]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[937]_i_3 
       (.I0(\f_permutation_l_/round_in [1512]),
        .I1(\f_permutation_l_/round_in [1447]),
        .I2(\out[1556]_i_8_n_0 ),
        .I3(\f_permutation_l_/round_in [1576]),
        .I4(\out[1556]_i_6_n_0 ),
        .O(\out[937]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[938]_i_1 
       (.I0(\f_permutation_l_/round_in [1124]),
        .I1(\out[1551]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[721] ),
        .I3(\out[1510]_i_3_n_0 ),
        .I4(\out[938]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [938]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[938]_i_2 
       (.I0(padder_out_1[92]),
        .I1(out[28]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1124]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[938]_i_3 
       (.I0(\f_permutation_l_/round_in [1513]),
        .I1(\f_permutation_l_/round_in [1448]),
        .I2(\out[1557]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1577]),
        .I4(\out[1557]_i_6_n_0 ),
        .O(\out[938]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[939]_i_1 
       (.I0(\f_permutation_l_/round_in [1125]),
        .I1(\out[1552]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[722] ),
        .I3(\out[1511]_i_3_n_0 ),
        .I4(\out[939]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [939]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[939]_i_2 
       (.I0(padder_out_1[93]),
        .I1(out[29]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1125]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[939]_i_3 
       (.I0(\f_permutation_l_/round_in [1514]),
        .I1(\f_permutation_l_/round_in [1449]),
        .I2(\out[1558]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1578]),
        .I4(\out[1558]_i_6_n_0 ),
        .O(\out[939]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[93]_i_1 
       (.I0(\out[1271]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[628] ),
        .I2(\f_permutation_l_/out_reg_n_0_[219] ),
        .I3(\out[1287]_i_3_n_0 ),
        .I4(\out[285]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [93]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[940]_i_1 
       (.I0(\f_permutation_l_/round_in [1126]),
        .I1(\out[1553]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[723] ),
        .I3(\out[1512]_i_3_n_0 ),
        .I4(\out[940]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [940]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[940]_i_2 
       (.I0(padder_out_1[94]),
        .I1(out[30]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1126]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[940]_i_3 
       (.I0(\f_permutation_l_/round_in [1515]),
        .I1(\f_permutation_l_/round_in [1450]),
        .I2(\out[1559]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1579]),
        .I4(\out[1559]_i_6_n_0 ),
        .O(\out[940]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[941]_i_1 
       (.I0(\f_permutation_l_/round_in [1127]),
        .I1(\out[1554]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[724] ),
        .I3(\out[1513]_i_3_n_0 ),
        .I4(\out[941]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [941]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[941]_i_2 
       (.I0(padder_out_1[95]),
        .I1(out[31]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1127]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[941]_i_3 
       (.I0(\f_permutation_l_/round_in [1516]),
        .I1(\f_permutation_l_/round_in [1451]),
        .I2(\out[1560]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1580]),
        .I4(\out[1560]_i_6_n_0 ),
        .O(\out[941]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[942]_i_1 
       (.I0(\f_permutation_l_/round_in [1128]),
        .I1(\out[1555]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[725] ),
        .I3(\out[1514]_i_3_n_0 ),
        .I4(\out[942]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [942]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[942]_i_2 
       (.I0(padder_out_1[80]),
        .I1(out[16]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1128]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[942]_i_3 
       (.I0(\f_permutation_l_/round_in [1517]),
        .I1(\f_permutation_l_/round_in [1452]),
        .I2(\out[1561]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1581]),
        .I4(\out[1561]_i_6_n_0 ),
        .O(\out[942]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF99F0660)) 
    \out[943]_i_1 
       (.I0(\f_permutation_l_/round_in [1129]),
        .I1(\out[1556]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[726] ),
        .I3(\out[1515]_i_3_n_0 ),
        .I4(\out[943]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [943]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[943]_i_2 
       (.I0(padder_out_1[81]),
        .I1(out[17]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1129]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[943]_i_3 
       (.I0(\f_permutation_l_/round_in [1518]),
        .I1(\f_permutation_l_/round_in [1453]),
        .I2(\out[1562]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1582]),
        .I4(\out[1562]_i_6_n_0 ),
        .O(\out[943]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[944]_i_1 
       (.I0(\f_permutation_l_/round_in [1130]),
        .I1(\out[1557]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[727] ),
        .I3(\out[1516]_i_3_n_0 ),
        .I4(\out[944]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [944]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[944]_i_2 
       (.I0(padder_out_1[82]),
        .I1(out[18]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1130]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[944]_i_3 
       (.I0(\f_permutation_l_/round_in [1519]),
        .I1(\f_permutation_l_/round_in [1454]),
        .I2(\out[1563]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1583]),
        .I4(\out[1563]_i_6_n_0 ),
        .O(\out[944]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[945]_i_1 
       (.I0(\f_permutation_l_/round_in [1131]),
        .I1(\out[1558]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[728] ),
        .I3(\out[1517]_i_3_n_0 ),
        .I4(\out[945]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [945]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[945]_i_2 
       (.I0(padder_out_1[83]),
        .I1(out[19]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1131]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[945]_i_3 
       (.I0(\f_permutation_l_/round_in [1520]),
        .I1(\f_permutation_l_/round_in [1455]),
        .I2(\out[1564]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1584]),
        .I4(\out[1564]_i_6_n_0 ),
        .O(\out[945]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[946]_i_1 
       (.I0(\f_permutation_l_/round_in [1132]),
        .I1(\out[1559]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[729] ),
        .I3(\out[1518]_i_3_n_0 ),
        .I4(\out[946]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [946]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[946]_i_2 
       (.I0(padder_out_1[84]),
        .I1(out[20]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1132]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[946]_i_3 
       (.I0(\f_permutation_l_/round_in [1521]),
        .I1(\f_permutation_l_/round_in [1456]),
        .I2(\out[1565]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1585]),
        .I4(\out[1565]_i_6_n_0 ),
        .O(\out[946]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[947]_i_1 
       (.I0(\f_permutation_l_/round_in [1133]),
        .I1(\out[1560]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[730] ),
        .I3(\out[1519]_i_3_n_0 ),
        .I4(\out[947]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [947]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[947]_i_2 
       (.I0(padder_out_1[85]),
        .I1(out[21]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1133]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[947]_i_3 
       (.I0(\f_permutation_l_/round_in [1522]),
        .I1(\f_permutation_l_/round_in [1457]),
        .I2(\out[1566]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1586]),
        .I4(\out[1566]_i_6_n_0 ),
        .O(\out[947]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[948]_i_1 
       (.I0(\f_permutation_l_/round_in [1134]),
        .I1(\out[1561]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[731] ),
        .I3(\out[1520]_i_3_n_0 ),
        .I4(\out[948]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [948]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[948]_i_2 
       (.I0(padder_out_1[86]),
        .I1(out[22]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1134]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[948]_i_3 
       (.I0(\f_permutation_l_/round_in [1523]),
        .I1(\f_permutation_l_/round_in [1458]),
        .I2(\out[1567]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1587]),
        .I4(\out[1567]_i_9_n_0 ),
        .O(\out[948]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[949]_i_1 
       (.I0(\f_permutation_l_/round_in [1135]),
        .I1(\out[1562]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[732] ),
        .I3(\out[1521]_i_3_n_0 ),
        .I4(\out[949]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [949]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[949]_i_2 
       (.I0(padder_out_1[87]),
        .I1(out[23]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1135]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[949]_i_3 
       (.I0(\f_permutation_l_/round_in [1524]),
        .I1(\f_permutation_l_/round_in [1459]),
        .I2(\out[1568]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1588]),
        .I4(\out[1568]_i_6_n_0 ),
        .O(\out[949]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[94]_i_1 
       (.I0(\out[1272]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[629] ),
        .I2(\f_permutation_l_/out_reg_n_0_[220] ),
        .I3(\out[1544]_i_3_n_0 ),
        .I4(\out[286]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [94]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[950]_i_1 
       (.I0(\f_permutation_l_/round_in [1136]),
        .I1(\out[1563]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[733] ),
        .I3(\out[1522]_i_3_n_0 ),
        .I4(\out[950]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [950]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[950]_i_2 
       (.I0(padder_out_1[72]),
        .I1(out[8]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1136]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[950]_i_3 
       (.I0(\f_permutation_l_/round_in [1525]),
        .I1(\f_permutation_l_/round_in [1460]),
        .I2(\out[1569]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1589]),
        .I4(\out[1569]_i_6_n_0 ),
        .O(\out[950]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[951]_i_1 
       (.I0(\f_permutation_l_/round_in [1137]),
        .I1(\out[1564]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[734] ),
        .I3(\out[1523]_i_3_n_0 ),
        .I4(\out[951]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [951]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[951]_i_2 
       (.I0(padder_out_1[73]),
        .I1(out[9]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1137]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[951]_i_3 
       (.I0(\f_permutation_l_/round_in [1526]),
        .I1(\f_permutation_l_/round_in [1461]),
        .I2(\out[1570]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1590]),
        .I4(\out[1570]_i_6_n_0 ),
        .O(\out[951]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[952]_i_1 
       (.I0(\f_permutation_l_/round_in [1138]),
        .I1(\out[1565]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[735] ),
        .I3(\out[1524]_i_3_n_0 ),
        .I4(\out[952]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [952]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[952]_i_2 
       (.I0(padder_out_1[74]),
        .I1(out[10]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1138]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[952]_i_3 
       (.I0(\f_permutation_l_/round_in [1527]),
        .I1(\f_permutation_l_/round_in [1462]),
        .I2(\out[1571]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1591]),
        .I4(\out[1571]_i_6_n_0 ),
        .O(\out[952]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[953]_i_1 
       (.I0(\f_permutation_l_/round_in [1139]),
        .I1(\out[1566]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[736] ),
        .I3(\out[1525]_i_3_n_0 ),
        .I4(\out[953]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [953]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[953]_i_2 
       (.I0(padder_out_1[75]),
        .I1(out[11]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1139]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[953]_i_3 
       (.I0(\f_permutation_l_/round_in [1528]),
        .I1(\f_permutation_l_/round_in [1463]),
        .I2(\out[1572]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1592]),
        .I4(\out[1572]_i_6_n_0 ),
        .O(\out[953]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[954]_i_1 
       (.I0(\f_permutation_l_/round_in [1140]),
        .I1(\out[1567]_i_3_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[737] ),
        .I3(\out[1526]_i_3_n_0 ),
        .I4(\out[954]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [954]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[954]_i_2 
       (.I0(padder_out_1[76]),
        .I1(out[12]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1140]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[954]_i_3 
       (.I0(\f_permutation_l_/round_in [1529]),
        .I1(\f_permutation_l_/round_in [1464]),
        .I2(\out[1573]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1593]),
        .I4(\out[1573]_i_6_n_0 ),
        .O(\out[954]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[955]_i_1 
       (.I0(\f_permutation_l_/round_in [1141]),
        .I1(\out[1568]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[738] ),
        .I3(\out[1527]_i_3_n_0 ),
        .I4(\out[955]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [955]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[955]_i_2 
       (.I0(padder_out_1[77]),
        .I1(out[13]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1141]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[955]_i_3 
       (.I0(\f_permutation_l_/round_in [1530]),
        .I1(\f_permutation_l_/round_in [1465]),
        .I2(\out[1574]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1594]),
        .I4(\out[1574]_i_6_n_0 ),
        .O(\out[955]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[956]_i_1 
       (.I0(\f_permutation_l_/round_in [1142]),
        .I1(\out[1569]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[739] ),
        .I3(\out[1528]_i_3_n_0 ),
        .I4(\out[956]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [956]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[956]_i_2 
       (.I0(padder_out_1[78]),
        .I1(out[14]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1142]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[956]_i_3 
       (.I0(\f_permutation_l_/round_in [1531]),
        .I1(\f_permutation_l_/round_in [1466]),
        .I2(\out[1575]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1595]),
        .I4(\out[1575]_i_6_n_0 ),
        .O(\out[956]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[957]_i_1 
       (.I0(\f_permutation_l_/round_in [1143]),
        .I1(\out[1570]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[740] ),
        .I3(\out[1529]_i_3_n_0 ),
        .I4(\out[957]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [957]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[957]_i_2 
       (.I0(padder_out_1[79]),
        .I1(out[15]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1143]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[957]_i_3 
       (.I0(\f_permutation_l_/round_in [1532]),
        .I1(\f_permutation_l_/round_in [1467]),
        .I2(\out[1576]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1596]),
        .I4(\out[1576]_i_6_n_0 ),
        .O(\out[957]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[958]_i_1 
       (.I0(\f_permutation_l_/round_in [1144]),
        .I1(\out[1571]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[741] ),
        .I3(\out[1530]_i_3_n_0 ),
        .I4(\out[958]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [958]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[958]_i_2 
       (.I0(padder_out_1[64]),
        .I1(out[0]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1144]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[958]_i_3 
       (.I0(\f_permutation_l_/round_in [1533]),
        .I1(\f_permutation_l_/round_in [1468]),
        .I2(\out[1577]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1597]),
        .I4(\out[1577]_i_6_n_0 ),
        .O(\out[958]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h9FF96006)) 
    \out[959]_i_1 
       (.I0(\f_permutation_l_/round_in [1145]),
        .I1(\out[1572]_i_4_n_0 ),
        .I2(\f_permutation_l_/out_reg_n_0_[742] ),
        .I3(\out[1531]_i_3_n_0 ),
        .I4(\out[959]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [959]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h6C)) 
    \out[959]_i_2 
       (.I0(padder_out_1[65]),
        .I1(out[1]),
        .I2(\out[1542]_i_6_n_0 ),
        .O(\f_permutation_l_/round_in [1145]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h96696996)) 
    \out[959]_i_3 
       (.I0(\f_permutation_l_/round_in [1534]),
        .I1(\f_permutation_l_/round_in [1469]),
        .I2(\out[1578]_i_7_n_0 ),
        .I3(\f_permutation_l_/round_in [1598]),
        .I4(\out[1578]_i_6_n_0 ),
        .O(\out[959]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[95]_i_1 
       (.I0(\out[1273]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[630] ),
        .I2(\f_permutation_l_/out_reg_n_0_[221] ),
        .I3(\out[1545]_i_3_n_0 ),
        .I4(\out[287]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [95]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[960]_i_1 
       (.I0(\out[1582]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[131] ),
        .I2(\out[1216]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1004] ),
        .I4(\out[1466]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [960]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[961]_i_1 
       (.I0(\out[1583]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[132] ),
        .I2(\out[1217]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1005] ),
        .I4(\out[1467]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [961]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[962]_i_1 
       (.I0(\out[1584]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[133] ),
        .I2(\out[1218]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1006] ),
        .I4(\out[1468]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [962]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[963]_i_1 
       (.I0(\out[1585]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[134] ),
        .I2(\out[1219]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1007] ),
        .I4(\out[1469]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [963]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[964]_i_1 
       (.I0(\out[1586]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[135] ),
        .I2(\out[1220]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1008] ),
        .I4(\out[1470]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [964]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[965]_i_1 
       (.I0(\out[1587]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[136] ),
        .I2(\out[1221]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1009] ),
        .I4(\out[1471]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [965]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[966]_i_1 
       (.I0(\out[1588]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[137] ),
        .I2(\out[1222]_i_2_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1010] ),
        .I4(\out[1408]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [966]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[967]_i_1 
       (.I0(\out[1589]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[138] ),
        .I2(\out[1223]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1011] ),
        .I4(\out[1409]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [967]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[968]_i_1 
       (.I0(\out[1590]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[139] ),
        .I2(\out[1224]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1012] ),
        .I4(\out[1410]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [968]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[969]_i_1 
       (.I0(\out[1591]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[140] ),
        .I2(\out[1225]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1013] ),
        .I4(\out[1411]_i_2_n_0 ),
        .O(\f_permutation_l_/round_out [969]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[96]_i_1 
       (.I0(\out[1274]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[631] ),
        .I2(\f_permutation_l_/out_reg_n_0_[222] ),
        .I3(\out[1546]_i_3_n_0 ),
        .I4(\out[288]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [96]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[970]_i_1 
       (.I0(\out[1592]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[141] ),
        .I2(\out[1226]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1014] ),
        .I4(\out[1412]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [970]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[971]_i_1 
       (.I0(\out[1593]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[142] ),
        .I2(\out[1227]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1015] ),
        .I4(\out[1413]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [971]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[972]_i_1 
       (.I0(\out[1594]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[143] ),
        .I2(\out[1228]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1016] ),
        .I4(\out[1414]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [972]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[973]_i_1 
       (.I0(\out[1595]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[144] ),
        .I2(\out[1229]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1017] ),
        .I4(\out[1415]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [973]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[974]_i_1 
       (.I0(\out[1596]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[145] ),
        .I2(\out[1230]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1018] ),
        .I4(\out[1416]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [974]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[975]_i_1 
       (.I0(\out[1597]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[146] ),
        .I2(\out[1231]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1019] ),
        .I4(\out[1417]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [975]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[976]_i_1 
       (.I0(\out[1598]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[147] ),
        .I2(\out[1232]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1020] ),
        .I4(\out[1418]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [976]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[977]_i_1 
       (.I0(\out[1599]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[148] ),
        .I2(\out[1233]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1021] ),
        .I4(\out[1419]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [977]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[978]_i_1 
       (.I0(\out[1472]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[149] ),
        .I2(\out[1234]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1022] ),
        .I4(\out[1420]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [978]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[979]_i_1 
       (.I0(\out[1537]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[150] ),
        .I2(\out[1235]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[1023] ),
        .I4(\out[1421]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [979]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[97]_i_1 
       (.I0(\out[1275]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[632] ),
        .I2(\f_permutation_l_/out_reg_n_0_[223] ),
        .I3(\out[1547]_i_3_n_0 ),
        .I4(\out[289]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [97]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[980]_i_1 
       (.I0(\out[1538]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[151] ),
        .I2(\out[1236]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[960] ),
        .I4(\out[1422]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [980]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h66696966)) 
    \out[981]_i_1 
       (.I0(\out[1045]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[152] ),
        .I2(\out[1237]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[961] ),
        .I4(\out[1423]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [981]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[982]_i_1 
       (.I0(\out[1540]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[153] ),
        .I2(\out[1238]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[962] ),
        .I4(\out[1424]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [982]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[983]_i_1 
       (.I0(\out[1541]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[154] ),
        .I2(\out[1239]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[963] ),
        .I4(\out[1425]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [983]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[984]_i_1 
       (.I0(\out[1542]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[155] ),
        .I2(\out[1240]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[964] ),
        .I4(\out[1426]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [984]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[985]_i_1 
       (.I0(\out[1543]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[156] ),
        .I2(\out[1241]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[965] ),
        .I4(\out[1427]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [985]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[986]_i_1 
       (.I0(\out[1544]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[157] ),
        .I2(\out[1242]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[966] ),
        .I4(\out[1428]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [986]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[987]_i_1 
       (.I0(\out[1545]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[158] ),
        .I2(\out[1243]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[967] ),
        .I4(\out[1429]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [987]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[988]_i_1 
       (.I0(\out[1546]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[159] ),
        .I2(\out[1244]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[968] ),
        .I4(\out[1430]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [988]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[989]_i_1 
       (.I0(\out[1547]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[160] ),
        .I2(\out[1245]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[969] ),
        .I4(\out[1431]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [989]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[98]_i_1 
       (.I0(\out[1276]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[633] ),
        .I2(\f_permutation_l_/out_reg_n_0_[224] ),
        .I3(\out[1548]_i_3_n_0 ),
        .I4(\out[290]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [98]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[990]_i_1 
       (.I0(\out[1548]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[161] ),
        .I2(\out[1246]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[970] ),
        .I4(\out[1432]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [990]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[991]_i_1 
       (.I0(\out[1549]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[162] ),
        .I2(\out[1247]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[971] ),
        .I4(\out[1433]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [991]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[992]_i_1 
       (.I0(\out[1550]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[163] ),
        .I2(\out[1248]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[972] ),
        .I4(\out[1434]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [992]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[993]_i_1 
       (.I0(\out[1551]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[164] ),
        .I2(\out[1249]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[973] ),
        .I4(\out[1435]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [993]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[994]_i_1 
       (.I0(\out[1552]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[165] ),
        .I2(\out[1250]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[974] ),
        .I4(\out[1436]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [994]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[995]_i_1 
       (.I0(\out[1553]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[166] ),
        .I2(\out[1251]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[975] ),
        .I4(\out[1437]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [995]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[996]_i_1 
       (.I0(\out[1554]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[167] ),
        .I2(\out[1252]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[976] ),
        .I4(\out[1438]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [996]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[997]_i_1 
       (.I0(\out[1555]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[168] ),
        .I2(\out[1253]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[977] ),
        .I4(\out[1439]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [997]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[998]_i_1 
       (.I0(\out[1556]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[169] ),
        .I2(\out[1254]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[978] ),
        .I4(\out[1440]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [998]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[999]_i_1 
       (.I0(\out[1557]_i_4_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[170] ),
        .I2(\out[1255]_i_3_n_0 ),
        .I3(\f_permutation_l_/out_reg_n_0_[979] ),
        .I4(\out[1441]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [999]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h69969999)) 
    \out[99]_i_1 
       (.I0(\out[1277]_i_2_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[634] ),
        .I2(\f_permutation_l_/out_reg_n_0_[225] ),
        .I3(\out[1549]_i_3_n_0 ),
        .I4(\out[291]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [99]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h99969699)) 
    \out[9]_i_1 
       (.I0(\out[1587]_i_3_n_0 ),
        .I1(\f_permutation_l_/out_reg_n_0_[199] ),
        .I2(\out[265]_i_3_n_0 ),
        .I3(\f_permutation_l_/round_in [1042]),
        .I4(\out[1511]_i_3_n_0 ),
        .O(\f_permutation_l_/round_out [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    out_ready_i_1
       (.I0(i),
        .I1(out_ready),
        .O(out_ready_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    out_ready_reg
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(out_ready_i_1_n_0),
        .Q(out_ready),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/done_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(done_i_1_n_0),
        .Q(\padder_l_/done ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[0] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[0]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[10] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[10]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[10] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[11] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[11]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[11] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[12] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[12]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[12] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[13] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[13]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[13] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[14] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[14]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[14] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[15] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[15]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[15] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[16] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[16]_i_1_n_0 ),
        .Q(\padder_l_/p_0_in ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[17] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[17]_i_1_n_0 ),
        .Q(buffer_full),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[1] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[1]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[2] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[2]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[3] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[3]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[4] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[4]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[5] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[5]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[6] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[6]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[7] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[7]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[7] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[8] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[8]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[8] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/i_reg[9] 
       (.C(clk),
        .CE(\padder_l_/i0 ),
        .D(\i[9]_i_1_n_0 ),
        .Q(\padder_l_/i_reg_n_0_[9] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF04)) 
    \padder_l_/out 
       (.I0(\padder_l_/done ),
        .I1(state),
        .I2(buffer_full),
        .I3(reset),
        .O(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'h88F0)) 
    \padder_l_/out[0]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[0]),
        .I3(is_last),
        .O(p_1_out[0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[10]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[10]),
        .I3(is_last),
        .O(p_1_out[10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[11]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[11]),
        .I3(is_last),
        .O(p_1_out[11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[12]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[12]),
        .I3(is_last),
        .O(p_1_out[12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[13]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[13]),
        .I3(is_last),
        .O(p_1_out[13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[14]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[14]),
        .I3(is_last),
        .O(p_1_out[14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[15]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[15]),
        .I3(is_last),
        .O(p_1_out[15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'hE2F0)) 
    \padder_l_/out[16]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[16]),
        .I3(is_last),
        .O(p_1_out[16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[17]_i_1 
       (.I0(byte_num[1]),
        .I1(in[17]),
        .I2(is_last),
        .O(p_1_out[17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[18]_i_1 
       (.I0(byte_num[1]),
        .I1(in[18]),
        .I2(is_last),
        .O(p_1_out[18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[19]_i_1 
       (.I0(byte_num[1]),
        .I1(in[19]),
        .I2(is_last),
        .O(p_1_out[19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[1]_i_1 
       (.I0(in[1]),
        .I1(is_last),
        .O(p_1_out[1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[20]_i_1 
       (.I0(byte_num[1]),
        .I1(in[20]),
        .I2(is_last),
        .O(p_1_out[20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[21]_i_1 
       (.I0(byte_num[1]),
        .I1(in[21]),
        .I2(is_last),
        .O(p_1_out[21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[22]_i_1 
       (.I0(byte_num[1]),
        .I1(in[22]),
        .I2(is_last),
        .O(p_1_out[22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT3 #(
    .INIT(8'h8C)) 
    \padder_l_/out[23]_i_1 
       (.I0(byte_num[1]),
        .I1(in[23]),
        .I2(is_last),
        .O(p_1_out[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'hF1F0)) 
    \padder_l_/out[24]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[24]),
        .I3(is_last),
        .O(p_1_out[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[25]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[25]),
        .I3(is_last),
        .O(p_1_out[25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[26]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[26]),
        .I3(is_last),
        .O(p_1_out[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[27]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[27]),
        .I3(is_last),
        .O(p_1_out[27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[28]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[28]),
        .I3(is_last),
        .O(p_1_out[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[29]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[29]),
        .I3(is_last),
        .O(p_1_out[29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[2]_i_1 
       (.I0(in[2]),
        .I1(is_last),
        .O(p_1_out[2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[30]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[30]),
        .I3(is_last),
        .O(p_1_out[30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'hE0F0)) 
    \padder_l_/out[31]_i_1 
       (.I0(byte_num[0]),
        .I1(byte_num[1]),
        .I2(in[31]),
        .I3(is_last),
        .O(p_1_out[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[3]_i_1 
       (.I0(in[3]),
        .I1(is_last),
        .O(p_1_out[3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[4]_i_1 
       (.I0(in[4]),
        .I1(is_last),
        .O(p_1_out[4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[5]_i_1 
       (.I0(in[5]),
        .I1(is_last),
        .O(p_1_out[5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \padder_l_/out[6]_i_1 
       (.I0(in[6]),
        .I1(is_last),
        .O(p_1_out[6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'hABA8)) 
    \padder_l_/out[7]_i_1 
       (.I0(\padder_l_/p_0_in ),
        .I1(state),
        .I2(is_last),
        .I3(in[7]),
        .O(p_1_out[7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'hA2F0)) 
    \padder_l_/out[8]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[8]),
        .I3(is_last),
        .O(p_1_out[8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'h80F0)) 
    \padder_l_/out[9]_i_1 
       (.I0(byte_num[1]),
        .I1(byte_num[0]),
        .I2(in[9]),
        .I3(is_last),
        .O(p_1_out[9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[0] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[0]),
        .Q(padder_out_1[0]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[100] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[68]),
        .Q(padder_out_1[100]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[101] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[69]),
        .Q(padder_out_1[101]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[102] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[70]),
        .Q(padder_out_1[102]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[103] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[71]),
        .Q(padder_out_1[103]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[104] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[72]),
        .Q(padder_out_1[104]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[105] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[73]),
        .Q(padder_out_1[105]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[106] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[74]),
        .Q(padder_out_1[106]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[107] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[75]),
        .Q(padder_out_1[107]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[108] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[76]),
        .Q(padder_out_1[108]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[109] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[77]),
        .Q(padder_out_1[109]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[10] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[10]),
        .Q(padder_out_1[10]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[110] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[78]),
        .Q(padder_out_1[110]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[111] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[79]),
        .Q(padder_out_1[111]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[112] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[80]),
        .Q(padder_out_1[112]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[113] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[81]),
        .Q(padder_out_1[113]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[114] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[82]),
        .Q(padder_out_1[114]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[115] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[83]),
        .Q(padder_out_1[115]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[116] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[84]),
        .Q(padder_out_1[116]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[117] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[85]),
        .Q(padder_out_1[117]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[118] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[86]),
        .Q(padder_out_1[118]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[119] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[87]),
        .Q(padder_out_1[119]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[11] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[11]),
        .Q(padder_out_1[11]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[120] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[88]),
        .Q(padder_out_1[120]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[121] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[89]),
        .Q(padder_out_1[121]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[122] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[90]),
        .Q(padder_out_1[122]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[123] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[91]),
        .Q(padder_out_1[123]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[124] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[92]),
        .Q(padder_out_1[124]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[125] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[93]),
        .Q(padder_out_1[125]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[126] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[94]),
        .Q(padder_out_1[126]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[127] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[95]),
        .Q(padder_out_1[127]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[128] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[96]),
        .Q(padder_out_1[128]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[129] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[97]),
        .Q(padder_out_1[129]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[12] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[12]),
        .Q(padder_out_1[12]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[130] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[98]),
        .Q(padder_out_1[130]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[131] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[99]),
        .Q(padder_out_1[131]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[132] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[100]),
        .Q(padder_out_1[132]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[133] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[101]),
        .Q(padder_out_1[133]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[134] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[102]),
        .Q(padder_out_1[134]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[135] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[103]),
        .Q(padder_out_1[135]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[136] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[104]),
        .Q(padder_out_1[136]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[137] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[105]),
        .Q(padder_out_1[137]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[138] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[106]),
        .Q(padder_out_1[138]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[139] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[107]),
        .Q(padder_out_1[139]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[13] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[13]),
        .Q(padder_out_1[13]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[140] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[108]),
        .Q(padder_out_1[140]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[141] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[109]),
        .Q(padder_out_1[141]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[142] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[110]),
        .Q(padder_out_1[142]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[143] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[111]),
        .Q(padder_out_1[143]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[144] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[112]),
        .Q(padder_out_1[144]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[145] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[113]),
        .Q(padder_out_1[145]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[146] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[114]),
        .Q(padder_out_1[146]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[147] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[115]),
        .Q(padder_out_1[147]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[148] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[116]),
        .Q(padder_out_1[148]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[149] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[117]),
        .Q(padder_out_1[149]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[14] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[14]),
        .Q(padder_out_1[14]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[150] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[118]),
        .Q(padder_out_1[150]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[151] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[119]),
        .Q(padder_out_1[151]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[152] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[120]),
        .Q(padder_out_1[152]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[153] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[121]),
        .Q(padder_out_1[153]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[154] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[122]),
        .Q(padder_out_1[154]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[155] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[123]),
        .Q(padder_out_1[155]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[156] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[124]),
        .Q(padder_out_1[156]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[157] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[125]),
        .Q(padder_out_1[157]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[158] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[126]),
        .Q(padder_out_1[158]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[159] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[127]),
        .Q(padder_out_1[159]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[15] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[15]),
        .Q(padder_out_1[15]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[160] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[128]),
        .Q(padder_out_1[160]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[161] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[129]),
        .Q(padder_out_1[161]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[162] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[130]),
        .Q(padder_out_1[162]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[163] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[131]),
        .Q(padder_out_1[163]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[164] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[132]),
        .Q(padder_out_1[164]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[165] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[133]),
        .Q(padder_out_1[165]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[166] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[134]),
        .Q(padder_out_1[166]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[167] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[135]),
        .Q(padder_out_1[167]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[168] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[136]),
        .Q(padder_out_1[168]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[169] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[137]),
        .Q(padder_out_1[169]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[16] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[16]),
        .Q(padder_out_1[16]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[170] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[138]),
        .Q(padder_out_1[170]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[171] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[139]),
        .Q(padder_out_1[171]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[172] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[140]),
        .Q(padder_out_1[172]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[173] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[141]),
        .Q(padder_out_1[173]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[174] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[142]),
        .Q(padder_out_1[174]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[175] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[143]),
        .Q(padder_out_1[175]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[176] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[144]),
        .Q(padder_out_1[176]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[177] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[145]),
        .Q(padder_out_1[177]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[178] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[146]),
        .Q(padder_out_1[178]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[179] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[147]),
        .Q(padder_out_1[179]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[17] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[17]),
        .Q(padder_out_1[17]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[180] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[148]),
        .Q(padder_out_1[180]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[181] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[149]),
        .Q(padder_out_1[181]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[182] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[150]),
        .Q(padder_out_1[182]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[183] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[151]),
        .Q(padder_out_1[183]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[184] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[152]),
        .Q(padder_out_1[184]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[185] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[153]),
        .Q(padder_out_1[185]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[186] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[154]),
        .Q(padder_out_1[186]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[187] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[155]),
        .Q(padder_out_1[187]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[188] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[156]),
        .Q(padder_out_1[188]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[189] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[157]),
        .Q(padder_out_1[189]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[18] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[18]),
        .Q(padder_out_1[18]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[190] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[158]),
        .Q(padder_out_1[190]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[191] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[159]),
        .Q(padder_out_1[191]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[192] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[160]),
        .Q(padder_out_1[192]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[193] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[161]),
        .Q(padder_out_1[193]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[194] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[162]),
        .Q(padder_out_1[194]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[195] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[163]),
        .Q(padder_out_1[195]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[196] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[164]),
        .Q(padder_out_1[196]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[197] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[165]),
        .Q(padder_out_1[197]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[198] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[166]),
        .Q(padder_out_1[198]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[199] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[167]),
        .Q(padder_out_1[199]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[19] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[19]),
        .Q(padder_out_1[19]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[1] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[1]),
        .Q(padder_out_1[1]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[200] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[168]),
        .Q(padder_out_1[200]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[201] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[169]),
        .Q(padder_out_1[201]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[202] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[170]),
        .Q(padder_out_1[202]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[203] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[171]),
        .Q(padder_out_1[203]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[204] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[172]),
        .Q(padder_out_1[204]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[205] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[173]),
        .Q(padder_out_1[205]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[206] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[174]),
        .Q(padder_out_1[206]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[207] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[175]),
        .Q(padder_out_1[207]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[208] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[176]),
        .Q(padder_out_1[208]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[209] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[177]),
        .Q(padder_out_1[209]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[20] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[20]),
        .Q(padder_out_1[20]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[210] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[178]),
        .Q(padder_out_1[210]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[211] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[179]),
        .Q(padder_out_1[211]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[212] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[180]),
        .Q(padder_out_1[212]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[213] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[181]),
        .Q(padder_out_1[213]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[214] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[182]),
        .Q(padder_out_1[214]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[215] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[183]),
        .Q(padder_out_1[215]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[216] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[184]),
        .Q(padder_out_1[216]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[217] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[185]),
        .Q(padder_out_1[217]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[218] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[186]),
        .Q(padder_out_1[218]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[219] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[187]),
        .Q(padder_out_1[219]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[21] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[21]),
        .Q(padder_out_1[21]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[220] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[188]),
        .Q(padder_out_1[220]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[221] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[189]),
        .Q(padder_out_1[221]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[222] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[190]),
        .Q(padder_out_1[222]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[223] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[191]),
        .Q(padder_out_1[223]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[224] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[192]),
        .Q(padder_out_1[224]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[225] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[193]),
        .Q(padder_out_1[225]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[226] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[194]),
        .Q(padder_out_1[226]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[227] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[195]),
        .Q(padder_out_1[227]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[228] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[196]),
        .Q(padder_out_1[228]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[229] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[197]),
        .Q(padder_out_1[229]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[22] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[22]),
        .Q(padder_out_1[22]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[230] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[198]),
        .Q(padder_out_1[230]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[231] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[199]),
        .Q(padder_out_1[231]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[232] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[200]),
        .Q(padder_out_1[232]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[233] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[201]),
        .Q(padder_out_1[233]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[234] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[202]),
        .Q(padder_out_1[234]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[235] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[203]),
        .Q(padder_out_1[235]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[236] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[204]),
        .Q(padder_out_1[236]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[237] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[205]),
        .Q(padder_out_1[237]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[238] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[206]),
        .Q(padder_out_1[238]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[239] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[207]),
        .Q(padder_out_1[239]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[23] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[23]),
        .Q(padder_out_1[23]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[240] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[208]),
        .Q(padder_out_1[240]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[241] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[209]),
        .Q(padder_out_1[241]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[242] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[210]),
        .Q(padder_out_1[242]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[243] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[211]),
        .Q(padder_out_1[243]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[244] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[212]),
        .Q(padder_out_1[244]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[245] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[213]),
        .Q(padder_out_1[245]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[246] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[214]),
        .Q(padder_out_1[246]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[247] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[215]),
        .Q(padder_out_1[247]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[248] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[216]),
        .Q(padder_out_1[248]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[249] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[217]),
        .Q(padder_out_1[249]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[24] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[24]),
        .Q(padder_out_1[24]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[250] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[218]),
        .Q(padder_out_1[250]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[251] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[219]),
        .Q(padder_out_1[251]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[252] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[220]),
        .Q(padder_out_1[252]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[253] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[221]),
        .Q(padder_out_1[253]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[254] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[222]),
        .Q(padder_out_1[254]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[255] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[223]),
        .Q(padder_out_1[255]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[256] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[224]),
        .Q(padder_out_1[256]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[257] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[225]),
        .Q(padder_out_1[257]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[258] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[226]),
        .Q(padder_out_1[258]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[259] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[227]),
        .Q(padder_out_1[259]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[25] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[25]),
        .Q(padder_out_1[25]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[260] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[228]),
        .Q(padder_out_1[260]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[261] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[229]),
        .Q(padder_out_1[261]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[262] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[230]),
        .Q(padder_out_1[262]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[263] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[231]),
        .Q(padder_out_1[263]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[264] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[232]),
        .Q(padder_out_1[264]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[265] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[233]),
        .Q(padder_out_1[265]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[266] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[234]),
        .Q(padder_out_1[266]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[267] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[235]),
        .Q(padder_out_1[267]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[268] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[236]),
        .Q(padder_out_1[268]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[269] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[237]),
        .Q(padder_out_1[269]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[26] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[26]),
        .Q(padder_out_1[26]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[270] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[238]),
        .Q(padder_out_1[270]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[271] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[239]),
        .Q(padder_out_1[271]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[272] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[240]),
        .Q(padder_out_1[272]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[273] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[241]),
        .Q(padder_out_1[273]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[274] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[242]),
        .Q(padder_out_1[274]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[275] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[243]),
        .Q(padder_out_1[275]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[276] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[244]),
        .Q(padder_out_1[276]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[277] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[245]),
        .Q(padder_out_1[277]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[278] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[246]),
        .Q(padder_out_1[278]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[279] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[247]),
        .Q(padder_out_1[279]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[27] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[27]),
        .Q(padder_out_1[27]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[280] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[248]),
        .Q(padder_out_1[280]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[281] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[249]),
        .Q(padder_out_1[281]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[282] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[250]),
        .Q(padder_out_1[282]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[283] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[251]),
        .Q(padder_out_1[283]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[284] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[252]),
        .Q(padder_out_1[284]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[285] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[253]),
        .Q(padder_out_1[285]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[286] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[254]),
        .Q(padder_out_1[286]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[287] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[255]),
        .Q(padder_out_1[287]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[288] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[256]),
        .Q(padder_out_1[288]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[289] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[257]),
        .Q(padder_out_1[289]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[28] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[28]),
        .Q(padder_out_1[28]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[290] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[258]),
        .Q(padder_out_1[290]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[291] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[259]),
        .Q(padder_out_1[291]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[292] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[260]),
        .Q(padder_out_1[292]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[293] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[261]),
        .Q(padder_out_1[293]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[294] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[262]),
        .Q(padder_out_1[294]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[295] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[263]),
        .Q(padder_out_1[295]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[296] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[264]),
        .Q(padder_out_1[296]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[297] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[265]),
        .Q(padder_out_1[297]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[298] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[266]),
        .Q(padder_out_1[298]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[299] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[267]),
        .Q(padder_out_1[299]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[29] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[29]),
        .Q(padder_out_1[29]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[2] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[2]),
        .Q(padder_out_1[2]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[300] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[268]),
        .Q(padder_out_1[300]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[301] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[269]),
        .Q(padder_out_1[301]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[302] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[270]),
        .Q(padder_out_1[302]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[303] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[271]),
        .Q(padder_out_1[303]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[304] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[272]),
        .Q(padder_out_1[304]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[305] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[273]),
        .Q(padder_out_1[305]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[306] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[274]),
        .Q(padder_out_1[306]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[307] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[275]),
        .Q(padder_out_1[307]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[308] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[276]),
        .Q(padder_out_1[308]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[309] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[277]),
        .Q(padder_out_1[309]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[30] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[30]),
        .Q(padder_out_1[30]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[310] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[278]),
        .Q(padder_out_1[310]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[311] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[279]),
        .Q(padder_out_1[311]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[312] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[280]),
        .Q(padder_out_1[312]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[313] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[281]),
        .Q(padder_out_1[313]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[314] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[282]),
        .Q(padder_out_1[314]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[315] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[283]),
        .Q(padder_out_1[315]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[316] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[284]),
        .Q(padder_out_1[316]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[317] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[285]),
        .Q(padder_out_1[317]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[318] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[286]),
        .Q(padder_out_1[318]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[319] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[287]),
        .Q(padder_out_1[319]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[31] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[31]),
        .Q(padder_out_1[31]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[320] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[288]),
        .Q(padder_out_1[320]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[321] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[289]),
        .Q(padder_out_1[321]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[322] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[290]),
        .Q(padder_out_1[322]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[323] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[291]),
        .Q(padder_out_1[323]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[324] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[292]),
        .Q(padder_out_1[324]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[325] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[293]),
        .Q(padder_out_1[325]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[326] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[294]),
        .Q(padder_out_1[326]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[327] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[295]),
        .Q(padder_out_1[327]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[328] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[296]),
        .Q(padder_out_1[328]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[329] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[297]),
        .Q(padder_out_1[329]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[32] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[0]),
        .Q(padder_out_1[32]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[330] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[298]),
        .Q(padder_out_1[330]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[331] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[299]),
        .Q(padder_out_1[331]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[332] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[300]),
        .Q(padder_out_1[332]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[333] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[301]),
        .Q(padder_out_1[333]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[334] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[302]),
        .Q(padder_out_1[334]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[335] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[303]),
        .Q(padder_out_1[335]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[336] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[304]),
        .Q(padder_out_1[336]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[337] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[305]),
        .Q(padder_out_1[337]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[338] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[306]),
        .Q(padder_out_1[338]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[339] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[307]),
        .Q(padder_out_1[339]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[33] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[1]),
        .Q(padder_out_1[33]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[340] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[308]),
        .Q(padder_out_1[340]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[341] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[309]),
        .Q(padder_out_1[341]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[342] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[310]),
        .Q(padder_out_1[342]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[343] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[311]),
        .Q(padder_out_1[343]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[344] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[312]),
        .Q(padder_out_1[344]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[345] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[313]),
        .Q(padder_out_1[345]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[346] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[314]),
        .Q(padder_out_1[346]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[347] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[315]),
        .Q(padder_out_1[347]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[348] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[316]),
        .Q(padder_out_1[348]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[349] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[317]),
        .Q(padder_out_1[349]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[34] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[2]),
        .Q(padder_out_1[34]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[350] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[318]),
        .Q(padder_out_1[350]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[351] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[319]),
        .Q(padder_out_1[351]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[352] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[320]),
        .Q(padder_out_1[352]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[353] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[321]),
        .Q(padder_out_1[353]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[354] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[322]),
        .Q(padder_out_1[354]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[355] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[323]),
        .Q(padder_out_1[355]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[356] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[324]),
        .Q(padder_out_1[356]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[357] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[325]),
        .Q(padder_out_1[357]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[358] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[326]),
        .Q(padder_out_1[358]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[359] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[327]),
        .Q(padder_out_1[359]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[35] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[3]),
        .Q(padder_out_1[35]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[360] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[328]),
        .Q(padder_out_1[360]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[361] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[329]),
        .Q(padder_out_1[361]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[362] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[330]),
        .Q(padder_out_1[362]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[363] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[331]),
        .Q(padder_out_1[363]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[364] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[332]),
        .Q(padder_out_1[364]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[365] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[333]),
        .Q(padder_out_1[365]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[366] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[334]),
        .Q(padder_out_1[366]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[367] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[335]),
        .Q(padder_out_1[367]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[368] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[336]),
        .Q(padder_out_1[368]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[369] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[337]),
        .Q(padder_out_1[369]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[36] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[4]),
        .Q(padder_out_1[36]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[370] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[338]),
        .Q(padder_out_1[370]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[371] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[339]),
        .Q(padder_out_1[371]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[372] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[340]),
        .Q(padder_out_1[372]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[373] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[341]),
        .Q(padder_out_1[373]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[374] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[342]),
        .Q(padder_out_1[374]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[375] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[343]),
        .Q(padder_out_1[375]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[376] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[344]),
        .Q(padder_out_1[376]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[377] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[345]),
        .Q(padder_out_1[377]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[378] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[346]),
        .Q(padder_out_1[378]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[379] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[347]),
        .Q(padder_out_1[379]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[37] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[5]),
        .Q(padder_out_1[37]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[380] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[348]),
        .Q(padder_out_1[380]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[381] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[349]),
        .Q(padder_out_1[381]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[382] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[350]),
        .Q(padder_out_1[382]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[383] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[351]),
        .Q(padder_out_1[383]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[384] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[352]),
        .Q(padder_out_1[384]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[385] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[353]),
        .Q(padder_out_1[385]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[386] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[354]),
        .Q(padder_out_1[386]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[387] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[355]),
        .Q(padder_out_1[387]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[388] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[356]),
        .Q(padder_out_1[388]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[389] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[357]),
        .Q(padder_out_1[389]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[38] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[6]),
        .Q(padder_out_1[38]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[390] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[358]),
        .Q(padder_out_1[390]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[391] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[359]),
        .Q(padder_out_1[391]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[392] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[360]),
        .Q(padder_out_1[392]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[393] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[361]),
        .Q(padder_out_1[393]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[394] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[362]),
        .Q(padder_out_1[394]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[395] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[363]),
        .Q(padder_out_1[395]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[396] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[364]),
        .Q(padder_out_1[396]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[397] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[365]),
        .Q(padder_out_1[397]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[398] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[366]),
        .Q(padder_out_1[398]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[399] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[367]),
        .Q(padder_out_1[399]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[39] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[7]),
        .Q(padder_out_1[39]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[3] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[3]),
        .Q(padder_out_1[3]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[400] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[368]),
        .Q(padder_out_1[400]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[401] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[369]),
        .Q(padder_out_1[401]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[402] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[370]),
        .Q(padder_out_1[402]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[403] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[371]),
        .Q(padder_out_1[403]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[404] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[372]),
        .Q(padder_out_1[404]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[405] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[373]),
        .Q(padder_out_1[405]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[406] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[374]),
        .Q(padder_out_1[406]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[407] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[375]),
        .Q(padder_out_1[407]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[408] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[376]),
        .Q(padder_out_1[408]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[409] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[377]),
        .Q(padder_out_1[409]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[40] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[8]),
        .Q(padder_out_1[40]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[410] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[378]),
        .Q(padder_out_1[410]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[411] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[379]),
        .Q(padder_out_1[411]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[412] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[380]),
        .Q(padder_out_1[412]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[413] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[381]),
        .Q(padder_out_1[413]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[414] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[382]),
        .Q(padder_out_1[414]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[415] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[383]),
        .Q(padder_out_1[415]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[416] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[384]),
        .Q(padder_out_1[416]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[417] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[385]),
        .Q(padder_out_1[417]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[418] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[386]),
        .Q(padder_out_1[418]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[419] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[387]),
        .Q(padder_out_1[419]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[41] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[9]),
        .Q(padder_out_1[41]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[420] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[388]),
        .Q(padder_out_1[420]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[421] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[389]),
        .Q(padder_out_1[421]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[422] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[390]),
        .Q(padder_out_1[422]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[423] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[391]),
        .Q(padder_out_1[423]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[424] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[392]),
        .Q(padder_out_1[424]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[425] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[393]),
        .Q(padder_out_1[425]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[426] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[394]),
        .Q(padder_out_1[426]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[427] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[395]),
        .Q(padder_out_1[427]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[428] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[396]),
        .Q(padder_out_1[428]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[429] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[397]),
        .Q(padder_out_1[429]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[42] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[10]),
        .Q(padder_out_1[42]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[430] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[398]),
        .Q(padder_out_1[430]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[431] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[399]),
        .Q(padder_out_1[431]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[432] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[400]),
        .Q(padder_out_1[432]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[433] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[401]),
        .Q(padder_out_1[433]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[434] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[402]),
        .Q(padder_out_1[434]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[435] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[403]),
        .Q(padder_out_1[435]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[436] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[404]),
        .Q(padder_out_1[436]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[437] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[405]),
        .Q(padder_out_1[437]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[438] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[406]),
        .Q(padder_out_1[438]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[439] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[407]),
        .Q(padder_out_1[439]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[43] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[11]),
        .Q(padder_out_1[43]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[440] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[408]),
        .Q(padder_out_1[440]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[441] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[409]),
        .Q(padder_out_1[441]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[442] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[410]),
        .Q(padder_out_1[442]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[443] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[411]),
        .Q(padder_out_1[443]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[444] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[412]),
        .Q(padder_out_1[444]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[445] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[413]),
        .Q(padder_out_1[445]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[446] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[414]),
        .Q(padder_out_1[446]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[447] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[415]),
        .Q(padder_out_1[447]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[448] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[416]),
        .Q(padder_out_1[448]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[449] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[417]),
        .Q(padder_out_1[449]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[44] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[12]),
        .Q(padder_out_1[44]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[450] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[418]),
        .Q(padder_out_1[450]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[451] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[419]),
        .Q(padder_out_1[451]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[452] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[420]),
        .Q(padder_out_1[452]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[453] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[421]),
        .Q(padder_out_1[453]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[454] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[422]),
        .Q(padder_out_1[454]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[455] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[423]),
        .Q(padder_out_1[455]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[456] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[424]),
        .Q(padder_out_1[456]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[457] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[425]),
        .Q(padder_out_1[457]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[458] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[426]),
        .Q(padder_out_1[458]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[459] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[427]),
        .Q(padder_out_1[459]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[45] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[13]),
        .Q(padder_out_1[45]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[460] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[428]),
        .Q(padder_out_1[460]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[461] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[429]),
        .Q(padder_out_1[461]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[462] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[430]),
        .Q(padder_out_1[462]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[463] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[431]),
        .Q(padder_out_1[463]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[464] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[432]),
        .Q(padder_out_1[464]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[465] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[433]),
        .Q(padder_out_1[465]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[466] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[434]),
        .Q(padder_out_1[466]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[467] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[435]),
        .Q(padder_out_1[467]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[468] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[436]),
        .Q(padder_out_1[468]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[469] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[437]),
        .Q(padder_out_1[469]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[46] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[14]),
        .Q(padder_out_1[46]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[470] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[438]),
        .Q(padder_out_1[470]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[471] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[439]),
        .Q(padder_out_1[471]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[472] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[440]),
        .Q(padder_out_1[472]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[473] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[441]),
        .Q(padder_out_1[473]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[474] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[442]),
        .Q(padder_out_1[474]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[475] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[443]),
        .Q(padder_out_1[475]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[476] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[444]),
        .Q(padder_out_1[476]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[477] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[445]),
        .Q(padder_out_1[477]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[478] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[446]),
        .Q(padder_out_1[478]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[479] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[447]),
        .Q(padder_out_1[479]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[47] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[15]),
        .Q(padder_out_1[47]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[480] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[448]),
        .Q(padder_out_1[480]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[481] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[449]),
        .Q(padder_out_1[481]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[482] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[450]),
        .Q(padder_out_1[482]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[483] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[451]),
        .Q(padder_out_1[483]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[484] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[452]),
        .Q(padder_out_1[484]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[485] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[453]),
        .Q(padder_out_1[485]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[486] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[454]),
        .Q(padder_out_1[486]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[487] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[455]),
        .Q(padder_out_1[487]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[488] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[456]),
        .Q(padder_out_1[488]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[489] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[457]),
        .Q(padder_out_1[489]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[48] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[16]),
        .Q(padder_out_1[48]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[490] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[458]),
        .Q(padder_out_1[490]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[491] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[459]),
        .Q(padder_out_1[491]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[492] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[460]),
        .Q(padder_out_1[492]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[493] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[461]),
        .Q(padder_out_1[493]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[494] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[462]),
        .Q(padder_out_1[494]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[495] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[463]),
        .Q(padder_out_1[495]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[496] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[464]),
        .Q(padder_out_1[496]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[497] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[465]),
        .Q(padder_out_1[497]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[498] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[466]),
        .Q(padder_out_1[498]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[499] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[467]),
        .Q(padder_out_1[499]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[49] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[17]),
        .Q(padder_out_1[49]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[4] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[4]),
        .Q(padder_out_1[4]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[500] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[468]),
        .Q(padder_out_1[500]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[501] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[469]),
        .Q(padder_out_1[501]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[502] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[470]),
        .Q(padder_out_1[502]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[503] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[471]),
        .Q(padder_out_1[503]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[504] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[472]),
        .Q(padder_out_1[504]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[505] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[473]),
        .Q(padder_out_1[505]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[506] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[474]),
        .Q(padder_out_1[506]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[507] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[475]),
        .Q(padder_out_1[507]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[508] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[476]),
        .Q(padder_out_1[508]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[509] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[477]),
        .Q(padder_out_1[509]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[50] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[18]),
        .Q(padder_out_1[50]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[510] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[478]),
        .Q(padder_out_1[510]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[511] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[479]),
        .Q(padder_out_1[511]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[512] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[480]),
        .Q(padder_out_1[512]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[513] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[481]),
        .Q(padder_out_1[513]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[514] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[482]),
        .Q(padder_out_1[514]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[515] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[483]),
        .Q(padder_out_1[515]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[516] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[484]),
        .Q(padder_out_1[516]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[517] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[485]),
        .Q(padder_out_1[517]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[518] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[486]),
        .Q(padder_out_1[518]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[519] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[487]),
        .Q(padder_out_1[519]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[51] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[19]),
        .Q(padder_out_1[51]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[520] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[488]),
        .Q(padder_out_1[520]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[521] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[489]),
        .Q(padder_out_1[521]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[522] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[490]),
        .Q(padder_out_1[522]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[523] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[491]),
        .Q(padder_out_1[523]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[524] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[492]),
        .Q(padder_out_1[524]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[525] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[493]),
        .Q(padder_out_1[525]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[526] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[494]),
        .Q(padder_out_1[526]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[527] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[495]),
        .Q(padder_out_1[527]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[528] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[496]),
        .Q(padder_out_1[528]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[529] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[497]),
        .Q(padder_out_1[529]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[52] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[20]),
        .Q(padder_out_1[52]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[530] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[498]),
        .Q(padder_out_1[530]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[531] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[499]),
        .Q(padder_out_1[531]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[532] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[500]),
        .Q(padder_out_1[532]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[533] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[501]),
        .Q(padder_out_1[533]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[534] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[502]),
        .Q(padder_out_1[534]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[535] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[503]),
        .Q(padder_out_1[535]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[536] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[504]),
        .Q(padder_out_1[536]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[537] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[505]),
        .Q(padder_out_1[537]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[538] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[506]),
        .Q(padder_out_1[538]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[539] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[507]),
        .Q(padder_out_1[539]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[53] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[21]),
        .Q(padder_out_1[53]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[540] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[508]),
        .Q(padder_out_1[540]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[541] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[509]),
        .Q(padder_out_1[541]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[542] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[510]),
        .Q(padder_out_1[542]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[543] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[511]),
        .Q(padder_out_1[543]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[544] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[512]),
        .Q(padder_out_1[544]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[545] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[513]),
        .Q(padder_out_1[545]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[546] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[514]),
        .Q(padder_out_1[546]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[547] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[515]),
        .Q(padder_out_1[547]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[548] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[516]),
        .Q(padder_out_1[548]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[549] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[517]),
        .Q(padder_out_1[549]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[54] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[22]),
        .Q(padder_out_1[54]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[550] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[518]),
        .Q(padder_out_1[550]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[551] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[519]),
        .Q(padder_out_1[551]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[552] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[520]),
        .Q(padder_out_1[552]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[553] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[521]),
        .Q(padder_out_1[553]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[554] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[522]),
        .Q(padder_out_1[554]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[555] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[523]),
        .Q(padder_out_1[555]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[556] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[524]),
        .Q(padder_out_1[556]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[557] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[525]),
        .Q(padder_out_1[557]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[558] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[526]),
        .Q(padder_out_1[558]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[559] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[527]),
        .Q(padder_out_1[559]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[55] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[23]),
        .Q(padder_out_1[55]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[560] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[528]),
        .Q(padder_out_1[560]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[561] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[529]),
        .Q(padder_out_1[561]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[562] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[530]),
        .Q(padder_out_1[562]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[563] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[531]),
        .Q(padder_out_1[563]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[564] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[532]),
        .Q(padder_out_1[564]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[565] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[533]),
        .Q(padder_out_1[565]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[566] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[534]),
        .Q(padder_out_1[566]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[567] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[535]),
        .Q(padder_out_1[567]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[568] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[536]),
        .Q(padder_out_1[568]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[569] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[537]),
        .Q(padder_out_1[569]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[56] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[24]),
        .Q(padder_out_1[56]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[570] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[538]),
        .Q(padder_out_1[570]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[571] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[539]),
        .Q(padder_out_1[571]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[572] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[540]),
        .Q(padder_out_1[572]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[573] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[541]),
        .Q(padder_out_1[573]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[574] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[542]),
        .Q(padder_out_1[574]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[575] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[543]),
        .Q(padder_out_1[575]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[57] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[25]),
        .Q(padder_out_1[57]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[58] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[26]),
        .Q(padder_out_1[58]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[59] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[27]),
        .Q(padder_out_1[59]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[5] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[5]),
        .Q(padder_out_1[5]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[60] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[28]),
        .Q(padder_out_1[60]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[61] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[29]),
        .Q(padder_out_1[61]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[62] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[30]),
        .Q(padder_out_1[62]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[63] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[31]),
        .Q(padder_out_1[63]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[64] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[32]),
        .Q(padder_out_1[64]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[65] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[33]),
        .Q(padder_out_1[65]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[66] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[34]),
        .Q(padder_out_1[66]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[67] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[35]),
        .Q(padder_out_1[67]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[68] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[36]),
        .Q(padder_out_1[68]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[69] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[37]),
        .Q(padder_out_1[69]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[6] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[6]),
        .Q(padder_out_1[6]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[70] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[38]),
        .Q(padder_out_1[70]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[71] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[39]),
        .Q(padder_out_1[71]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[72] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[40]),
        .Q(padder_out_1[72]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[73] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[41]),
        .Q(padder_out_1[73]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[74] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[42]),
        .Q(padder_out_1[74]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[75] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[43]),
        .Q(padder_out_1[75]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[76] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[44]),
        .Q(padder_out_1[76]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[77] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[45]),
        .Q(padder_out_1[77]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[78] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[46]),
        .Q(padder_out_1[78]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[79] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[47]),
        .Q(padder_out_1[79]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[7] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[7]),
        .Q(padder_out_1[7]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[80] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[48]),
        .Q(padder_out_1[80]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[81] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[49]),
        .Q(padder_out_1[81]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[82] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[50]),
        .Q(padder_out_1[82]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[83] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[51]),
        .Q(padder_out_1[83]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[84] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[52]),
        .Q(padder_out_1[84]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[85] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[53]),
        .Q(padder_out_1[85]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[86] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[54]),
        .Q(padder_out_1[86]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[87] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[55]),
        .Q(padder_out_1[87]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[88] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[56]),
        .Q(padder_out_1[88]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[89] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[57]),
        .Q(padder_out_1[89]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[8] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[8]),
        .Q(padder_out_1[8]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[90] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[58]),
        .Q(padder_out_1[90]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[91] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[59]),
        .Q(padder_out_1[91]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[92] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[60]),
        .Q(padder_out_1[92]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[93] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[61]),
        .Q(padder_out_1[93]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[94] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[62]),
        .Q(padder_out_1[94]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[95] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[63]),
        .Q(padder_out_1[95]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[96] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[64]),
        .Q(padder_out_1[96]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[97] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[65]),
        .Q(padder_out_1[97]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[98] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[66]),
        .Q(padder_out_1[98]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[99] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(padder_out_1[67]),
        .Q(padder_out_1[99]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/out_reg[9] 
       (.C(clk),
        .CE(\padder_l_/update__1 ),
        .D(p_1_out[9]),
        .Q(padder_out_1[9]),
        .R(\padder_l_/out_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \padder_l_/state_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(state_i_1_n_0),
        .Q(state),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0054)) 
    \padder_l_/update 
       (.I0(\padder_l_/done ),
        .I1(state),
        .I2(in_ready),
        .I3(buffer_full),
        .O(\padder_l_/update__1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF0054)) 
    \padder_l_/update__0 
       (.I0(\padder_l_/done ),
        .I1(state),
        .I2(in_ready),
        .I3(buffer_full),
        .I4(update__0_i_1_n_0),
        .O(\padder_l_/i0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT2 #(
    .INIT(4'hE)) 
    state_i_1
       (.I0(is_last),
        .I1(state),
        .O(state_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    update__0_i_1
       (.I0(buffer_full),
        .I1(\f_permutation_l_/calc ),
        .O(update__0_i_1_n_0));
endmodule
