module dfadd
   (clk,
    reset,
    start,
    finish,
    waitrequest,
    return_val);
  input clk;
  input reset;
  input start;
  output finish;
  input waitrequest;
  output [31:0]return_val;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_cur_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[2]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state[4]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire FSM_sequential_cur_state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_29_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_29_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_29_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_34_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_34_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_34_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_39_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_39_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_39_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_51_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_51_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_51_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_56_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_56_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_56_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_5_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_5_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_5_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_61_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_61_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_61_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_66_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_66_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_66_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_71_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_71_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_71_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_76_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_76_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_76_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_81_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_81_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_81_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_86_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_86_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_86_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_91_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_91_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[2]_i_91_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_34_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_34_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_34_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \FSM_sequential_cur_state_reg[4]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_15;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_17;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_19;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_24;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_25;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_27;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_28;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ONE_8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_136;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_137;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_138;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_139;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_140;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_142;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_143;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_144;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_145;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_146;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_147;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_148;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_149;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_150;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_151;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_152;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_153;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_154;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_155;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_156;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_157;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_158;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_159;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_160;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_161;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_162;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_163;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_164;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_165;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_166;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_167;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_168;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_169;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_170;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_171;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_172;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_173;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_174;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_175;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_176;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_177;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_178;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_227;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_228;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_234;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_237;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_245;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ZERO_249;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cur_state;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_100_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[1]_rep_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[2]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[4]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[5]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state[6]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire cur_state_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_22_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_22_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_22_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_29_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_29_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_29_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_34_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_34_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_34_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_43_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_43_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_43_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_48_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_48_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_48_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_55_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_55_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_61_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_61_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_61_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_72_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_72_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_72_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_73_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_73_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_73_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_85_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_85_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_85_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_90_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_90_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_90_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_94_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_94_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[1]_i_94_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_23_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_23_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_23_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_27_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_27_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_27_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_32_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_32_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[2]_i_32_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_15_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_15_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_15_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_16_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_29_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_29_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_29_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_38_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_38_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_38_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_43_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_43_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_43_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_52_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_52_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_52_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_65_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_65_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_65_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_74_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_74_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_74_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[5]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_18_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_18_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_18_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_20_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_20_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_20_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \cur_state_reg[6]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire finish;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire finish_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_101_zExp1ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_101_zExp1ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[11]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[11]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[11]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[11]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[15]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[19]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[23]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[27]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[31]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[31]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[31]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[31]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[3]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zExp1ii_reg_reg[7]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_101_zSig0i12i_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[12]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[16]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[20]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[24]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[28]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[32]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[36]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[40]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[44]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[44]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[44]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[63]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_101_zSig0i12i_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[16]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[20]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[24]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[28]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[32]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[36]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[40]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[44]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[44]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[44]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[44]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[60]_i_1_GND_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[63]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[63]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[63]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_101_zSig0i12i_reg_reg[63]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_103_105_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_121_aExp0ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_121_bExp0ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_136_expDiff0ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_136_expDiff0ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_158_159_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_159_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_158_160_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_158_160_reg[62]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_158_bExp1ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_169_expDiff1ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_191_192_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_191_193_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_191_193_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_191_aExp1ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_0ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_12_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_12_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_12_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_1_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_1_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_1_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_2_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_2_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_2_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_7_n_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_7_n_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_197_reg_reg_i_7_n_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_199_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_iiiii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_iiiii_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_195_zSig0ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[27]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[35]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[39]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[43]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[43]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[43]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[43]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[63]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[63]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_195_zSig0ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[19]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[19]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[19]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[23]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[23]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[23]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[27]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[27]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[27]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[31]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[31]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[31]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[35]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[35]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[35]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[39]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[39]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[39]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[43]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[43]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[43]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[43]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[47]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[47]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[47]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[47]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[51]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[51]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[51]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[51]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[55]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[55]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[55]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[55]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[59]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[59]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[59]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_195_zSig0ii_reg_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_1_2_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_2_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_2_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_1_4_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_1_main_result02_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_1_main_result02_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[0]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[0]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[0]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[0]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[12]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[16]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[20]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[24]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[28]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[28]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[28]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[28]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[4]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_main_result02_reg_reg[8]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_1_scevgep_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_1_scevgep_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[25]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[29]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[29]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[29]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[31]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_1_scevgep_reg_reg[31]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_27_expDiff0i2i_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_0i_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[10]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[11]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[12]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[13]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[14]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[17]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[18]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[1]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[20]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[21]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[22]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[24]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[25]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[26]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[28]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[29]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[30]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[32]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[34]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[38]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[40]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[41]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[42]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[42]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[42]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[43]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[43]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[43]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[44]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[44]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[44]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[45]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[45]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[46]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[46]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[46]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[47]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[47]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[47]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[48]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[48]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[48]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[49]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[50]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[50]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[50]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[51]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[51]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[51]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[51]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[51]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[52]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[52]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[52]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[52]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[53]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[54]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[54]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[54]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[55]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[55]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[55]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[56]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[56]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[56]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[58]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[58]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[58]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[59]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[59]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[5]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[60]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[60]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[60]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[61]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[61]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[61]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[62]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[7]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_float64_addexit_0i_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[15]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[15]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[15]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[19]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[19]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[19]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[23]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[23]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[23]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[32]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[3]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[3]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[3]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[3]_i_7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[62]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[7]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[7]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_0i_reg_reg[7]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_218_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg[3]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_float64_addexit_218_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[19]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[19]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[19]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[23]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[23]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[23]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[27]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[27]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[27]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_14_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_14_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_14_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_24_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_24_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_24_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[3]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_218_reg_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_220_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_float64_addexit_220_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[16]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[16]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[16]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[20]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[20]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[20]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[24]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[24]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[24]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[28]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[28]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[28]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[31]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[4]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[4]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[4]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_float64_addexit_220_reg_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_float64_addexit_exitcond1_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:0]\main_inst/A ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [42:1]\main_inst/C ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/CI ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg[6]_rep_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/cur_state_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:23]\main_inst/data2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/data24 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [32:0]\main_inst/data5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/finish_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_102_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zExp1ii1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_101_zExp1ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_101_zSig0i12i_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_103_105_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_103_107 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_103_107_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_112_114 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_121_122 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_121_aExp0ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_121_bExp0ii_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_123_124 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_127_128 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_136_139_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:1]\main_inst/main_136_141_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:0]\main_inst/main_136_expDiff0ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_145_152 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_154_156 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_158_159 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:0]\main_inst/main_158_159_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_158_160 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [62:10]\main_inst/main_158_160_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_158_bExp1ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_158_bExp1ii_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:9]\main_inst/main_15_17 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_15_17_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:9]\main_inst/main_15_19_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_165_166 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_169_172_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_169_expDiff1ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_175_176 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_177_185 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_187_189 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_191_192 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [62:10]\main_inst/main_191_192_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_191_193 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:0]\main_inst/main_191_193_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_191_aExp1ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_191_aExp1ii_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_0ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_195_196 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]\main_inst/main_195_196_reg_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg[31]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg[8]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg[8]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg[8]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_196_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_197 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_197_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_199 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:24]\main_inst/main_195_200 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:24]\main_inst/main_195_200_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:24]\main_inst/main_195_asinkiiii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:24]\main_inst/main_195_extracttiiii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_iiiii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_iiiii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zExp0ii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zExp0ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/main_195_zSig0ii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_2_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_2_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_2_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_2_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_3_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_1_main_result02_reg_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:23]\main_inst/main_1_scevgep ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:3]\main_inst/main_1_scevgep_reg1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_1_scevgep_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_23_24 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_27_30_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_27_expDiff0i2i_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_33_34 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_35_43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_35_44 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_45_47 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_59_62_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [5:1]\main_inst/main_59_64_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [0:0]\main_inst/main_59_expDiff1i3i_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_68_75 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_68_76 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_81_83 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:9]\main_inst/main_91_92 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_0i121_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_0i129_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_0i13_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [62:0]\main_inst/main_float64_addexit_0i_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_0i_reg0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_0i_reg_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_float64_addexit_218 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_218_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/main_float64_addexit_220 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_220_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_exitcond1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_float64_addexit_exitcond1_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_shift64RightJammingexit3ii_z0i2ii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:0]\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_shift64RightJammingexit9ii_94_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:40]\main_inst/main_shift64RightJammingexit9ii_95 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [40:0]\main_inst/main_shift64RightJammingexit9ii_95_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/main_shift64RightJammingexit9ii_99_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [62:1]\main_inst/main_shift64RightJammingexit9ii_ii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:10]\main_inst/main_shift64RightJammingexitii_z0iii ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [41:0]\main_inst/main_shift64RightJammingexitii_z0iii_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [6:0]\main_inst/next_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [4:0]\main_inst/roundAndPackFloat64/cur_state ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/return_val_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_11_16_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_19_20 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_21_29 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_31_33 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_4_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_6_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:63]\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_35 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:11]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:52]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:52]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:10]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:1]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_39 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [9:0]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:8]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:8]\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_57_0_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/roundAndPackFloat64_arg_zExp ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/roundAndPackFloat64_arg_zSig ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSign ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_arg_zSign_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_finish ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_finish_reg1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_finish_reg_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_memory_controller_enable_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\main_inst/roundAndPackFloat64_memory_controller_in_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_memory_controller_write_enable_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [63:0]\main_inst/roundAndPackFloat64_return_val_reg ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_start ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_inst/roundAndPackFloat64_start_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_normalizeRoundAndPackFloat64exitii_209_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_209_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_209_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexit3ii_z0i2ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_shift64RightJammingexit3ii_z0i2ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexit9ii_100_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_100_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexit9ii_94_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[0]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[16]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[34]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[34]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[36]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[38]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[38]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[40]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[6]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_shift64RightJammingexit9ii_94_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexit9ii_95_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_106_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_119_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_120_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_121_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_122_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_123_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_124_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_125_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_126_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_127_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_128_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_129_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_130_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_131_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_132_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_133_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_135_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_136_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_137_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_140_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_145_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_146_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_147_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_148_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_149_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_150_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_151_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_152_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_153_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_154_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_155_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_156_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_157_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_158_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_159_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_160_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_161_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_162_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_163_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_164_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_165_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_166_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_167_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_168_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_169_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_170_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_171_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_172_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_173_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_174_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_175_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_178_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_179_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_180_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_181_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_182_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_183_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_184_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_185_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_186_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_187_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_188_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_189_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_190_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_191_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_192_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_193_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_194_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_195_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_196_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_197_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_198_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_199_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_200_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_201_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_202_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_203_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_204_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_205_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_206_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_207_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_208_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_209_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_210_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_211_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_212_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_213_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_215_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_216_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[16]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[33]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[34]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[35]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[36]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[37]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[38]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_shift64RightJammingexit9ii_95_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexit9ii_ii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[11]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[11]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[11]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[15]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[15]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[19]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[19]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[19]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[23]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[23]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[23]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[27]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[27]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[27]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[27]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[35]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[35]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[35]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[35]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[39]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[39]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[39]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[39]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[43]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[43]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[43]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[43]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[48]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[7]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[7]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[7]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg[7]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_shift64RightJammingexit9ii_ii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[48]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[48]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[63]_i_1_VCC_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire main_shift64RightJammingexitii_z0iii_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_119_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_120_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_121_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_122_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_123_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_124_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_125_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_126_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_127_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_128_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_129_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_132_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_133_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_136_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_137_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_140_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_145_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_146_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_147_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_148_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_149_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_150_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_151_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_152_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_153_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_154_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_155_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_156_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_157_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_158_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_159_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_160_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_161_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_162_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_163_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_164_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_165_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_166_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_167_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_168_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_169_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_170_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_171_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_172_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_173_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_176_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_177_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_178_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_179_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_180_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_181_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_182_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_183_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_184_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_185_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_186_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_187_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_188_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_189_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_190_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_191_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_192_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_193_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_194_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_195_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_196_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_197_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_198_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_199_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_200_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_201_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_202_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_203_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_205_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_206_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_207_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_208_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_209_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_210_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[41]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[41]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[8]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[9]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]main_shift64RightJammingexitii_z0iii_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:23]memory_controller_address_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_address_b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_enable_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_enable_b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_enable_reg_a_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_enable_reg_a_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_enable_reg_b_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire memory_controller_in_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\memory_controller_inst/float_exception_flags/q_a_wire ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\memory_controller_inst/float_exception_flags/q_b_wire ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/float_exception_flags/ram_reg_ENBWREN_cooolgate_en_sig_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/float_exception_flags_write_enable_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/memory_controller_enable_reg_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/memory_controller_enable_reg_b ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\memory_controller_inst/memory_controller_out_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]\memory_controller_inst/memory_controller_out_b ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/select_float_exception_flags_reg_a ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \memory_controller_inst/select_float_exception_flags_reg_b ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]memory_controller_out_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]memory_controller_out_b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_47_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_48_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_49_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_50_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_51_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_52_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_53_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_54_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_55_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_56_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_57_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_58_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_59_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_60_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_61_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_63_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_64_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_65_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_66_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_67_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire ram_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire reset;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [31:0]return_val;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \return_val[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_11_16_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_11_16_reg[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_57_0_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[55]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[59]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[59]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[59]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[59]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]roundAndPackFloat64_57_0_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_arg_zExp;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[11]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[11]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[11]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[15]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[19]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[23]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[27]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[31]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[3]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[3]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[7]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[7]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[7]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]roundAndPackFloat64_arg_zExp_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_arg_zSig;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[2]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[31]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[32]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[33]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[34]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[35]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[36]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[37]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[38]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[40]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[41]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[42]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[42]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[43]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[43]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[43]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[44]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[44]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[44]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[45]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[45]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[45]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[46]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[46]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[46]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[47]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[47]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[47]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[47]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[48]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[48]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[48]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[48]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[49]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[49]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[49]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[4]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[50]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[50]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[50]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[50]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[51]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[51]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[51]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[51]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[52]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[52]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[52]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[52]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[53]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[53]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[53]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[54]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[54]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[54]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[54]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[55]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[55]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[55]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[56]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[56]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[56]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[57]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[58]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[58]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[58]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[59]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[5]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[60]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[61]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[62]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[63]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[6]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[7]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]roundAndPackFloat64_arg_zSig_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_arg_zSign;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_arg_zSign[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_finish_reg_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_return_val_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_return_val_reg[63]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_return_val_reg[63]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_shift64RightJammingexit_z0i_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_101_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_102_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_103_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_107_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_108_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_109_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_110_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_112_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_113_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_114_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_115_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_116_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_117_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_120_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_121_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_122_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_123_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_124_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_125_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_126_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_127_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_128_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_129_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_132_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_133_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_134_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_135_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_136_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_137_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_138_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_139_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_140_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_146_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_147_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_148_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_149_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_150_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_151_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_152_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_153_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_154_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_155_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_158_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_159_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_160_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_163_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_164_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_165_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_166_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_168_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_169_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_170_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_171_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_172_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_173_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_174_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_175_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_179_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_181_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_182_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_183_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_184_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_185_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_186_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_187_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_188_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_189_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_190_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_191_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_192_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_193_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_194_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_195_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_196_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_197_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_198_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_199_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_200_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_201_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_202_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_204_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_205_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_206_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_207_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_208_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_209_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_210_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_211_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_212_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_213_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_214_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_215_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_216_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_217_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_218_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_219_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_220_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_221_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_222_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_223_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_224_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_225_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_226_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_227_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_228_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_229_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_48_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_49_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_51_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_53_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_54_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_56_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_58_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_60_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_62_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_64_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_65_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_66_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_67_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_69_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_70_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_71_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_72_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_74_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_75_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_76_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_77_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_78_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_79_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_82_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_83_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_84_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_87_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_92_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_93_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_94_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_95_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_99_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_start_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_start_i_2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_start_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_start_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_50_reg_i_9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_55_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg[0]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]roundAndPackFloat64_thread6_55_reg_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread6_roundBits09_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread6_roundBits09_reg[9]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread_02_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[10]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[11]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_02_reg[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire roundAndPackFloat64_thread_roundBits0_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \roundAndPackFloat64_thread_roundBits0_reg[9]_i_6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire select_float_exception_flags_reg_a;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]select_float_exception_flags_reg_a_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_16_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_16_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_16_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_16_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_9_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_a_reg[1]_i_9_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire select_float_exception_flags_reg_b;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b[1]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b[1]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b[1]_i_4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b[1]_i_5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [3:0]select_float_exception_flags_reg_b_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_3 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_4 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_5 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_6 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \select_float_exception_flags_reg_b_reg[1]_i_8_n_7 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire start;

  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \FSM_sequential_cur_state[0]_i_1 
       (.I0(\FSM_sequential_cur_state[0]_i_2_n_0 ),
        .I1(\FSM_sequential_cur_state[0]_i_3_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I3(\FSM_sequential_cur_state[0]_i_4_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I5(\FSM_sequential_cur_state[0]_i_5_n_0 ),
        .O(FSM_sequential_cur_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00CD)) 
    \FSM_sequential_cur_state[0]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .O(\FSM_sequential_cur_state[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFC44)) 
    \FSM_sequential_cur_state[0]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_19_20 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [2]),
        .O(\FSM_sequential_cur_state[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h400C400F)) 
    \FSM_sequential_cur_state[0]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_6_7 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_3 ),
        .O(\FSM_sequential_cur_state[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFDF)) 
    \FSM_sequential_cur_state[0]_i_5 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_4_5 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .O(\FSM_sequential_cur_state[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    \FSM_sequential_cur_state[0]_i_6 
       (.I0(\FSM_sequential_cur_state[4]_i_10_n_0 ),
        .I1(\FSM_sequential_cur_state[0]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I5(\FSM_sequential_cur_state[4]_i_12_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_3 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[0]_i_7 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\FSM_sequential_cur_state[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h1167AAAA)) 
    \FSM_sequential_cur_state[1]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_4_5 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .O(\FSM_sequential_cur_state[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h033303000C1C0C1C)) 
    \FSM_sequential_cur_state[1]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_19_20 ),
        .I5(\main_inst/roundAndPackFloat64/cur_state [1]),
        .O(\FSM_sequential_cur_state[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_cur_state[2]_i_14 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .O(\FSM_sequential_cur_state[2]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_15 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ),
        .O(\FSM_sequential_cur_state[2]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_16 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ),
        .O(\FSM_sequential_cur_state[2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_17 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ),
        .O(\FSM_sequential_cur_state[2]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_18 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ),
        .O(\FSM_sequential_cur_state[2]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h03FFCB00)) 
    \FSM_sequential_cur_state[2]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_39 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [2]),
        .O(\FSM_sequential_cur_state[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_25 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ),
        .O(\FSM_sequential_cur_state[2]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_26 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ),
        .O(\FSM_sequential_cur_state[2]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_27 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ),
        .O(\FSM_sequential_cur_state[2]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_28 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ),
        .O(\FSM_sequential_cur_state[2]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3333FFFFECEF2020)) 
    \FSM_sequential_cur_state[2]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_19_20 ),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [2]),
        .O(\FSM_sequential_cur_state[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_35 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ),
        .O(\FSM_sequential_cur_state[2]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_36 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ),
        .O(\FSM_sequential_cur_state[2]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_37 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ),
        .O(\FSM_sequential_cur_state[2]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_38 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ),
        .O(\FSM_sequential_cur_state[2]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \FSM_sequential_cur_state[2]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[8] ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[2] ),
        .I4(\FSM_sequential_cur_state[2]_i_7_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_39 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[2]_i_44 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .O(\FSM_sequential_cur_state[2]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[2]_i_45 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\FSM_sequential_cur_state[2]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[2]_i_46 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\FSM_sequential_cur_state[2]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[2]_i_47 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ),
        .O(\FSM_sequential_cur_state[2]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[2]_i_48 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\FSM_sequential_cur_state[2]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[2]_i_49 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\FSM_sequential_cur_state[2]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[2]_i_50 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\FSM_sequential_cur_state[2]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_sequential_cur_state[2]_i_7 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[7] ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[9] ),
        .O(\FSM_sequential_cur_state[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \FSM_sequential_cur_state[2]_i_98 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .O(\FSM_sequential_cur_state[2]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB38C8C80BC8C8C80)) 
    \FSM_sequential_cur_state[3]_i_1 
       (.I0(\FSM_sequential_cur_state[3]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [4]),
        .O(\FSM_sequential_cur_state[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000FFFEE)) 
    \FSM_sequential_cur_state[3]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_35 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [2]),
        .O(\FSM_sequential_cur_state[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h555FFFFF555FFFFE)) 
    \FSM_sequential_cur_state[4]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I5(\main_inst/roundAndPackFloat64_start_reg_n_0 ),
        .O(\FSM_sequential_cur_state[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \FSM_sequential_cur_state[4]_i_10 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ),
        .O(\FSM_sequential_cur_state[4]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_sequential_cur_state[4]_i_11 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ),
        .O(\FSM_sequential_cur_state[4]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000000000000000)) 
    \FSM_sequential_cur_state[4]_i_12 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ),
        .O(\FSM_sequential_cur_state[4]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_cur_state[4]_i_14 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .O(\FSM_sequential_cur_state[4]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_15 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ),
        .O(\FSM_sequential_cur_state[4]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_16 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ),
        .O(\FSM_sequential_cur_state[4]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_17 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ),
        .O(\FSM_sequential_cur_state[4]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_18 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ),
        .O(\FSM_sequential_cur_state[4]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_19 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ),
        .O(\FSM_sequential_cur_state[4]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hC800FFFFC8000000)) 
    \FSM_sequential_cur_state[4]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_35 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I5(\FSM_sequential_cur_state[4]_i_4_n_0 ),
        .O(\FSM_sequential_cur_state[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_20 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ),
        .O(\FSM_sequential_cur_state[4]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_21 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ),
        .O(\FSM_sequential_cur_state[4]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_22 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ),
        .O(\FSM_sequential_cur_state[4]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_23 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ),
        .O(\FSM_sequential_cur_state[4]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_24 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ),
        .O(\FSM_sequential_cur_state[4]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_26 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ),
        .O(\FSM_sequential_cur_state[4]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_27 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ),
        .O(\FSM_sequential_cur_state[4]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_28 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ),
        .O(\FSM_sequential_cur_state[4]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_29 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ),
        .O(\FSM_sequential_cur_state[4]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \FSM_sequential_cur_state[4]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [1]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [8]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [3]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [5]),
        .I4(\FSM_sequential_cur_state[4]_i_5_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_35 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_30 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ),
        .O(\FSM_sequential_cur_state[4]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_31 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ),
        .O(\FSM_sequential_cur_state[4]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_32 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ),
        .O(\FSM_sequential_cur_state[4]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_33 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ),
        .O(\FSM_sequential_cur_state[4]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_35 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ),
        .O(\FSM_sequential_cur_state[4]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \FSM_sequential_cur_state[4]_i_36 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ),
        .O(\FSM_sequential_cur_state[4]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_37 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ),
        .O(\FSM_sequential_cur_state[4]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \FSM_sequential_cur_state[4]_i_38 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ),
        .O(\FSM_sequential_cur_state[4]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_cur_state[4]_i_39 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ),
        .O(\FSM_sequential_cur_state[4]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFBFF3F30000C0F0)) 
    \FSM_sequential_cur_state[4]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_6_7 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_4_5 ),
        .I4(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [4]),
        .O(\FSM_sequential_cur_state[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[4]_i_40 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ),
        .O(\FSM_sequential_cur_state[4]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[4]_i_41 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ),
        .O(\FSM_sequential_cur_state[4]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[4]_i_42 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\FSM_sequential_cur_state[4]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \FSM_sequential_cur_state[4]_i_43 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\FSM_sequential_cur_state[4]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \FSM_sequential_cur_state[4]_i_44 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\FSM_sequential_cur_state[4]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \FSM_sequential_cur_state[4]_i_5 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [9]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [0]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [4]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [6]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [2]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [7]),
        .O(\FSM_sequential_cur_state[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00040000)) 
    \FSM_sequential_cur_state[4]_i_6 
       (.I0(\FSM_sequential_cur_state[4]_i_8_n_0 ),
        .I1(\FSM_sequential_cur_state[4]_i_9_n_0 ),
        .I2(\FSM_sequential_cur_state[4]_i_10_n_0 ),
        .I3(\FSM_sequential_cur_state[4]_i_11_n_0 ),
        .I4(\FSM_sequential_cur_state[4]_i_12_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_6_7 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF7FFFFFFF)) 
    \FSM_sequential_cur_state[4]_i_8 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\FSM_sequential_cur_state[4]_i_22_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\FSM_sequential_cur_state[4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \FSM_sequential_cur_state[4]_i_9 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ),
        .I4(\FSM_sequential_cur_state[4]_i_23_n_0 ),
        .I5(\FSM_sequential_cur_state[4]_i_24_n_0 ),
        .O(\FSM_sequential_cur_state[4]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_cur_state_reg[1]_i_1 
       (.I0(\FSM_sequential_cur_state[1]_i_2_n_0 ),
        .I1(\FSM_sequential_cur_state[1]_i_3_n_0 ),
        .O(FSM_sequential_cur_state_reg),
        .S(\main_inst/roundAndPackFloat64/cur_state [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \FSM_sequential_cur_state_reg[2]_i_1 
       (.I0(\FSM_sequential_cur_state[2]_i_2_n_0 ),
        .I1(\FSM_sequential_cur_state[2]_i_3_n_0 ),
        .O(\FSM_sequential_cur_state_reg[2]_i_1_n_0 ),
        .S(\main_inst/roundAndPackFloat64/cur_state [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_13 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_24_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_13_n_0 ,\FSM_sequential_cur_state_reg[2]_i_13_n_1 ,\FSM_sequential_cur_state_reg[2]_i_13_n_2 ,\FSM_sequential_cur_state_reg[2]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\FSM_sequential_cur_state[2]_i_25_n_0 ,\FSM_sequential_cur_state[2]_i_26_n_0 ,\FSM_sequential_cur_state[2]_i_27_n_0 ,\FSM_sequential_cur_state[2]_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_19 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_29_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_19_n_0 ,\FSM_sequential_cur_state_reg[2]_i_19_n_1 ,\FSM_sequential_cur_state_reg[2]_i_19_n_2 ,\FSM_sequential_cur_state_reg[2]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_24 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_34_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_24_n_0 ,\FSM_sequential_cur_state_reg[2]_i_24_n_1 ,\FSM_sequential_cur_state_reg[2]_i_24_n_2 ,\FSM_sequential_cur_state_reg[2]_i_24_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\FSM_sequential_cur_state[2]_i_35_n_0 ,\FSM_sequential_cur_state[2]_i_36_n_0 ,\FSM_sequential_cur_state[2]_i_37_n_0 ,\FSM_sequential_cur_state[2]_i_38_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_29 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_39_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_29_n_0 ,\FSM_sequential_cur_state_reg[2]_i_29_n_1 ,\FSM_sequential_cur_state_reg[2]_i_29_n_2 ,\FSM_sequential_cur_state_reg[2]_i_29_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_34 
       (.CI(\<const0>__0__0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_34_n_0 ,\FSM_sequential_cur_state_reg[2]_i_34_n_1 ,\FSM_sequential_cur_state_reg[2]_i_34_n_2 ,\FSM_sequential_cur_state_reg[2]_i_34_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\FSM_sequential_cur_state[2]_i_44_n_0 ,\FSM_sequential_cur_state[2]_i_45_n_0 ,\FSM_sequential_cur_state[2]_i_46_n_0 }),
        .S({\FSM_sequential_cur_state[2]_i_47_n_0 ,\FSM_sequential_cur_state[2]_i_48_n_0 ,\FSM_sequential_cur_state[2]_i_49_n_0 ,\FSM_sequential_cur_state[2]_i_50_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_39 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_51_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_39_n_0 ,\FSM_sequential_cur_state_reg[2]_i_39_n_1 ,\FSM_sequential_cur_state_reg[2]_i_39_n_2 ,\FSM_sequential_cur_state_reg[2]_i_39_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_5 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_8_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ,\FSM_sequential_cur_state_reg[2]_i_5_n_5 ,\FSM_sequential_cur_state_reg[2]_i_5_n_6 ,\FSM_sequential_cur_state_reg[2]_i_5_n_7 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_51 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_56_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_51_n_0 ,\FSM_sequential_cur_state_reg[2]_i_51_n_1 ,\FSM_sequential_cur_state_reg[2]_i_51_n_2 ,\FSM_sequential_cur_state_reg[2]_i_51_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_56 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_61_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_56_n_0 ,\FSM_sequential_cur_state_reg[2]_i_56_n_1 ,\FSM_sequential_cur_state_reg[2]_i_56_n_2 ,\FSM_sequential_cur_state_reg[2]_i_56_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_6 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_13_n_0 ),
        .CO({\main_inst/roundAndPackFloat64/roundAndPackFloat64_19_20 ,\FSM_sequential_cur_state_reg[2]_i_6_n_1 ,\FSM_sequential_cur_state_reg[2]_i_6_n_2 ,\FSM_sequential_cur_state_reg[2]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\FSM_sequential_cur_state[2]_i_14_n_0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\FSM_sequential_cur_state[2]_i_15_n_0 ,\FSM_sequential_cur_state[2]_i_16_n_0 ,\FSM_sequential_cur_state[2]_i_17_n_0 ,\FSM_sequential_cur_state[2]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_61 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_66_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_61_n_0 ,\FSM_sequential_cur_state_reg[2]_i_61_n_1 ,\FSM_sequential_cur_state_reg[2]_i_61_n_2 ,\FSM_sequential_cur_state_reg[2]_i_61_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_66 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_71_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_66_n_0 ,\FSM_sequential_cur_state_reg[2]_i_66_n_1 ,\FSM_sequential_cur_state_reg[2]_i_66_n_2 ,\FSM_sequential_cur_state_reg[2]_i_66_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_71 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_76_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_71_n_0 ,\FSM_sequential_cur_state_reg[2]_i_71_n_1 ,\FSM_sequential_cur_state_reg[2]_i_71_n_2 ,\FSM_sequential_cur_state_reg[2]_i_71_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_76 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_81_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_76_n_0 ,\FSM_sequential_cur_state_reg[2]_i_76_n_1 ,\FSM_sequential_cur_state_reg[2]_i_76_n_2 ,\FSM_sequential_cur_state_reg[2]_i_76_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_8 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_19_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_8_n_0 ,\FSM_sequential_cur_state_reg[2]_i_8_n_1 ,\FSM_sequential_cur_state_reg[2]_i_8_n_2 ,\FSM_sequential_cur_state_reg[2]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_81 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_86_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_81_n_0 ,\FSM_sequential_cur_state_reg[2]_i_81_n_1 ,\FSM_sequential_cur_state_reg[2]_i_81_n_2 ,\FSM_sequential_cur_state_reg[2]_i_81_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_86 
       (.CI(\FSM_sequential_cur_state_reg[2]_i_91_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_86_n_0 ,\FSM_sequential_cur_state_reg[2]_i_86_n_1 ,\FSM_sequential_cur_state_reg[2]_i_86_n_2 ,\FSM_sequential_cur_state_reg[2]_i_86_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[2]_i_91 
       (.CI(\<const0>__0__0 ),
        .CO({\FSM_sequential_cur_state_reg[2]_i_91_n_0 ,\FSM_sequential_cur_state_reg[2]_i_91_n_1 ,\FSM_sequential_cur_state_reg[2]_i_91_n_2 ,\FSM_sequential_cur_state_reg[2]_i_91_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ,\<const0>__0__0 }),
        .S({\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ,\FSM_sequential_cur_state[2]_i_98_n_0 ,\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[4]_i_13 
       (.CI(\FSM_sequential_cur_state_reg[4]_i_25_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[4]_i_13_n_0 ,\FSM_sequential_cur_state_reg[4]_i_13_n_1 ,\FSM_sequential_cur_state_reg[4]_i_13_n_2 ,\FSM_sequential_cur_state_reg[4]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\FSM_sequential_cur_state[4]_i_26_n_0 ,\FSM_sequential_cur_state[4]_i_27_n_0 ,\FSM_sequential_cur_state[4]_i_28_n_0 ,\FSM_sequential_cur_state[4]_i_29_n_0 }),
        .S({\FSM_sequential_cur_state[4]_i_30_n_0 ,\FSM_sequential_cur_state[4]_i_31_n_0 ,\FSM_sequential_cur_state[4]_i_32_n_0 ,\FSM_sequential_cur_state[4]_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[4]_i_25 
       (.CI(\FSM_sequential_cur_state_reg[4]_i_34_n_0 ),
        .CO({\FSM_sequential_cur_state_reg[4]_i_25_n_0 ,\FSM_sequential_cur_state_reg[4]_i_25_n_1 ,\FSM_sequential_cur_state_reg[4]_i_25_n_2 ,\FSM_sequential_cur_state_reg[4]_i_25_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\FSM_sequential_cur_state[4]_i_35_n_0 ,\FSM_sequential_cur_state[4]_i_36_n_0 ,\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ,\<const0>__0__0 }),
        .S({\FSM_sequential_cur_state[4]_i_37_n_0 ,\FSM_sequential_cur_state[4]_i_38_n_0 ,\FSM_sequential_cur_state[4]_i_39_n_0 ,\FSM_sequential_cur_state[4]_i_40_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[4]_i_34 
       (.CI(\<const0>__0__0 ),
        .CO({\FSM_sequential_cur_state_reg[4]_i_34_n_0 ,\FSM_sequential_cur_state_reg[4]_i_34_n_1 ,\FSM_sequential_cur_state_reg[4]_i_34_n_2 ,\FSM_sequential_cur_state_reg[4]_i_34_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] }),
        .S({\FSM_sequential_cur_state[4]_i_41_n_0 ,\FSM_sequential_cur_state[4]_i_42_n_0 ,\FSM_sequential_cur_state[4]_i_43_n_0 ,\FSM_sequential_cur_state[4]_i_44_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \FSM_sequential_cur_state_reg[4]_i_7 
       (.CI(\FSM_sequential_cur_state_reg[4]_i_13_n_0 ),
        .CO({\main_inst/roundAndPackFloat64/roundAndPackFloat64_4_5 ,\FSM_sequential_cur_state_reg[4]_i_7_n_1 ,\FSM_sequential_cur_state_reg[4]_i_7_n_2 ,\FSM_sequential_cur_state_reg[4]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\FSM_sequential_cur_state[4]_i_14_n_0 ,\FSM_sequential_cur_state[4]_i_15_n_0 ,\FSM_sequential_cur_state[4]_i_16_n_0 ,\FSM_sequential_cur_state[4]_i_17_n_0 }),
        .S({\FSM_sequential_cur_state[4]_i_18_n_0 ,\FSM_sequential_cur_state[4]_i_19_n_0 ,\FSM_sequential_cur_state[4]_i_20_n_0 ,\FSM_sequential_cur_state[4]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_140
       (.G(ZERO_136));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_141
       (.G(ZERO_137));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_142
       (.G(ZERO_138));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_143
       (.G(ZERO_139));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_144
       (.G(ZERO_140));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_146
       (.G(ZERO_142));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_147
       (.G(ZERO_143));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_148
       (.G(ZERO_144));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_149
       (.G(ZERO_145));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_150
       (.G(ZERO_146));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_151
       (.G(ZERO_147));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_152
       (.G(ZERO_148));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_153
       (.G(ZERO_149));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_154
       (.G(ZERO_150));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_155
       (.G(ZERO_151));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_156
       (.G(ZERO_152));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_157
       (.G(ZERO_153));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_158
       (.G(ZERO_154));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_159
       (.G(ZERO_155));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_160
       (.G(ZERO_156));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_161
       (.G(ZERO_157));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_162
       (.G(ZERO_158));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_163
       (.G(ZERO_159));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_164
       (.G(ZERO_160));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_165
       (.G(ZERO_161));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_166
       (.G(ZERO_162));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_167
       (.G(ZERO_163));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_168
       (.G(ZERO_164));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_169
       (.G(ZERO_165));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_170
       (.G(ZERO_166));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_171
       (.G(ZERO_167));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_172
       (.G(ZERO_168));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_173
       (.G(ZERO_169));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_174
       (.G(ZERO_170));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_175
       (.G(ZERO_171));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_176
       (.G(ZERO_172));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_177
       (.G(ZERO_173));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_178
       (.G(ZERO_174));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_179
       (.G(ZERO_175));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_180
       (.G(ZERO_176));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_181
       (.G(ZERO_177));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_182
       (.G(ZERO_178));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_231
       (.G(ZERO_227));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_232
       (.G(ZERO_228));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_238
       (.G(ZERO_234));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_241
       (.G(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_249
       (.G(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND_253
       (.G(ZERO_249));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_53
       (.P(ONE_7));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_54
       (.P(ONE_8));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_56
       (.P(ONE_10));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_57
       (.P(ONE_11));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_58
       (.P(ONE_12));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_59
       (.P(ONE_13));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_60
       (.P(ONE_14));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_61
       (.P(ONE_15));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_62
       (.P(ONE_16));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_63
       (.P(ONE_17));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_64
       (.P(ONE_18));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_65
       (.P(ONE_19));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_66
       (.P(ONE_20));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_67
       (.P(ONE_21));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_68
       (.P(ONE_22));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_69
       (.P(ONE_23));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_70
       (.P(ONE_24));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_71
       (.P(ONE_25));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_73
       (.P(ONE_27));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC_74
       (.P(ONE_28));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \cur_state[0]_i_1 
       (.I0(\cur_state[0]_i_2_n_0 ),
        .I1(\cur_state[0]_i_3_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\cur_state_reg[0]_i_4_n_0 ),
        .I4(\cur_state[1]_i_5_n_0 ),
        .I5(\cur_state_reg[0]_i_5_n_0 ),
        .O(\main_inst/next_state [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2E0C22F0EEFF2EFF)) 
    \cur_state[0]_i_10 
       (.I0(cur_state_reg),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(cur_state));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h2F)) 
    \cur_state[0]_i_11 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h50003FFF)) 
    \cur_state[0]_i_12 
       (.I0(\main_inst/main_123_124 ),
        .I1(\main_inst/main_121_122 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \cur_state[0]_i_13 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h707F)) 
    \cur_state[0]_i_14 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCB)) 
    \cur_state[0]_i_16 
       (.I0(\main_inst/main_33_34 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \cur_state[0]_i_17 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFFFFFF4000)) 
    \cur_state[0]_i_2 
       (.I0(\cur_state[1]_i_7_n_0 ),
        .I1(\cur_state[1]_i_8_n_0 ),
        .I2(\cur_state[1]_i_9_n_0 ),
        .I3(\cur_state[1]_i_10_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h40FFFFFF40FF0000)) 
    \cur_state[0]_i_3 
       (.I0(\main_inst/main_float64_addexit_exitcond1_reg ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\cur_state[0]_i_6_n_0 ),
        .O(\cur_state[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h83BF83BC)) 
    \cur_state[0]_i_6 
       (.I0(\cur_state[3]_i_5_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/main_175_176 ),
        .O(\cur_state[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBF)) 
    \cur_state[0]_i_9 
       (.I0(\cur_state[6]_i_13_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \cur_state[1]_i_1 
       (.I0(\cur_state[1]_i_2_n_0 ),
        .I1(\cur_state[1]_i_3_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\cur_state[1]_i_4_n_0 ),
        .I4(\cur_state[1]_i_5_n_0 ),
        .I5(\cur_state_reg[1]_i_6_n_0 ),
        .O(\main_inst/next_state [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \cur_state[1]_i_10 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_ ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[4] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[6] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[7] ),
        .I4(\cur_state[1]_i_21_n_0 ),
        .O(\cur_state[1]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_100 
       (.I0(\main_inst/main_15_19_reg [17]),
        .I1(\main_inst/main_15_19_reg [16]),
        .I2(\main_inst/main_15_19_reg [15]),
        .O(\cur_state[1]_i_100_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_101 
       (.I0(\main_inst/main_15_19_reg [14]),
        .I1(\main_inst/main_15_19_reg [13]),
        .I2(\main_inst/main_15_19_reg [12]),
        .O(\cur_state[1]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_102 
       (.I0(\main_inst/main_15_19_reg [11]),
        .I1(\main_inst/main_15_19_reg [10]),
        .I2(\main_inst/main_15_19_reg [9]),
        .O(\cur_state[1]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h70)) 
    \cur_state[1]_i_12 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h08F80BF8)) 
    \cur_state[1]_i_13 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/main_127_128 ),
        .O(\cur_state[1]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hA0FF3F00)) 
    \cur_state[1]_i_14 
       (.I0(\main_inst/main_123_124 ),
        .I1(\main_inst/main_121_122 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0340)) 
    \cur_state[1]_i_15 
       (.I0(\main_inst/main_112_114 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4F000000)) 
    \cur_state[1]_i_16 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[1]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFAFACCFC0A0ACC0C)) 
    \cur_state[1]_i_17 
       (.I0(\cur_state_reg[1]_i_26_n_0 ),
        .I1(\cur_state[1]_i_27_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\cur_state[1]_i_28_n_0 ),
        .O(\cur_state[1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \cur_state[1]_i_18 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[20] ),
        .O(\cur_state[1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cur_state[1]_i_19 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[24] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[27] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[26] ),
        .O(\cur_state[1]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000FFFFFFFFBFFF)) 
    \cur_state[1]_i_2 
       (.I0(\cur_state[1]_i_7_n_0 ),
        .I1(\cur_state[1]_i_8_n_0 ),
        .I2(\cur_state[1]_i_9_n_0 ),
        .I3(\cur_state[1]_i_10_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \cur_state[1]_i_20 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[9] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[8] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[10] ),
        .O(\cur_state[1]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \cur_state[1]_i_21 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[2] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[1] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[5] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[3] ),
        .O(\cur_state[1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_23 
       (.I0(\main_inst/main_169_expDiff1ii_reg [30]),
        .I1(\main_inst/main_169_expDiff1ii_reg [31]),
        .O(\cur_state[1]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0370)) 
    \cur_state[1]_i_27 
       (.I0(\main_inst/main_23_24 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h38)) 
    \cur_state[1]_i_28 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h40FFEF0040FFEF05)) 
    \cur_state[1]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\cur_state[3]_i_5_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_inst/main_175_176 ),
        .O(\cur_state[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_30 
       (.I0(\main_inst/main_169_expDiff1ii_reg [28]),
        .I1(\main_inst/main_169_expDiff1ii_reg [29]),
        .O(\cur_state[1]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_31 
       (.I0(\main_inst/main_169_expDiff1ii_reg [26]),
        .I1(\main_inst/main_169_expDiff1ii_reg [27]),
        .O(\cur_state[1]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_32 
       (.I0(\main_inst/main_169_expDiff1ii_reg [24]),
        .I1(\main_inst/main_169_expDiff1ii_reg [25]),
        .O(\cur_state[1]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_33 
       (.I0(\main_inst/main_169_expDiff1ii_reg [22]),
        .I1(\main_inst/main_169_expDiff1ii_reg [23]),
        .O(\cur_state[1]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \cur_state[1]_i_4 
       (.I0(\cur_state[1]_i_12_n_0 ),
        .I1(\cur_state[1]_i_13_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\cur_state[1]_i_14_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\cur_state[1]_i_15_n_0 ),
        .O(\cur_state[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h38)) 
    \cur_state[1]_i_41 
       (.I0(\main_inst/main_33_34 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hBC)) 
    \cur_state[1]_i_42 
       (.I0(\main_inst/data24 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[1]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_44 
       (.I0(\main_inst/main_169_expDiff1ii_reg [20]),
        .I1(\main_inst/main_169_expDiff1ii_reg [21]),
        .O(\cur_state[1]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_45 
       (.I0(\main_inst/main_169_expDiff1ii_reg [18]),
        .I1(\main_inst/main_169_expDiff1ii_reg [19]),
        .O(\cur_state[1]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_46 
       (.I0(\main_inst/main_169_expDiff1ii_reg [16]),
        .I1(\main_inst/main_169_expDiff1ii_reg [17]),
        .O(\cur_state[1]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_47 
       (.I0(\main_inst/main_169_expDiff1ii_reg [14]),
        .I1(\main_inst/main_169_expDiff1ii_reg [15]),
        .O(\cur_state[1]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \cur_state[1]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .O(\cur_state[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_56 
       (.I0(\main_inst/main_169_expDiff1ii_reg [6]),
        .I1(\main_inst/main_169_expDiff1ii_reg [7]),
        .O(\cur_state[1]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_57 
       (.I0(\main_inst/main_169_expDiff1ii_reg [12]),
        .I1(\main_inst/main_169_expDiff1ii_reg [13]),
        .O(\cur_state[1]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_58 
       (.I0(\main_inst/main_169_expDiff1ii_reg [10]),
        .I1(\main_inst/main_169_expDiff1ii_reg [11]),
        .O(\cur_state[1]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_59 
       (.I0(\main_inst/main_169_expDiff1ii_reg [8]),
        .I1(\main_inst/main_169_expDiff1ii_reg [9]),
        .O(\cur_state[1]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \cur_state[1]_i_60 
       (.I0(\main_inst/main_169_expDiff1ii_reg [6]),
        .I1(\main_inst/main_169_expDiff1ii_reg [7]),
        .O(\cur_state[1]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_62 
       (.I0(\main_inst/main_103_107_reg [41]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .I2(\main_inst/main_103_107_reg [40]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .I5(\main_inst/main_103_107_reg [39]),
        .O(\cur_state[1]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_63 
       (.I0(\main_inst/main_103_107_reg [38]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I2(\main_inst/main_103_107_reg [37]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I5(\main_inst/main_103_107_reg [36]),
        .O(\cur_state[1]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_64 
       (.I0(\main_inst/main_103_107_reg [35]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_103_107_reg [34]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .I5(\main_inst/main_103_107_reg [33]),
        .O(\cur_state[1]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    \cur_state[1]_i_7 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[17] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[19] ),
        .I4(\cur_state[1]_i_18_n_0 ),
        .O(\cur_state[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_74 
       (.I0(\main_inst/main_103_107_reg [32]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I2(\main_inst/main_103_107_reg [31]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I5(\main_inst/main_103_107_reg [30]),
        .O(\cur_state[1]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_75 
       (.I0(\main_inst/main_103_107_reg [29]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .I2(\main_inst/main_103_107_reg [28]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .I5(\main_inst/main_103_107_reg [27]),
        .O(\cur_state[1]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_76 
       (.I0(\main_inst/main_103_107_reg [26]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_103_107_reg [25]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I5(\main_inst/main_103_107_reg [24]),
        .O(\cur_state[1]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_77 
       (.I0(\main_inst/main_103_107_reg [23]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .I2(\main_inst/main_103_107_reg [22]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .I5(\main_inst/main_103_107_reg [21]),
        .O(\cur_state[1]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \cur_state[1]_i_8 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[29] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[31] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[30] ),
        .I4(\cur_state[1]_i_19_n_0 ),
        .O(\cur_state[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_86 
       (.I0(\main_inst/main_103_107_reg [20]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_103_107_reg [19]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I5(\main_inst/main_103_107_reg [18]),
        .O(\cur_state[1]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_87 
       (.I0(\main_inst/main_103_107_reg [17]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .I2(\main_inst/main_103_107_reg [16]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .I5(\main_inst/main_103_107_reg [15]),
        .O(\cur_state[1]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[1]_i_88 
       (.I0(\main_inst/main_103_107_reg [14]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_103_107_reg [13]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .I4(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I5(\main_inst/main_103_107_reg [12]),
        .O(\cur_state[1]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \cur_state[1]_i_89 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I1(\main_inst/main_103_107_reg [10]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_103_107_reg [11]),
        .O(\cur_state[1]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \cur_state[1]_i_9 
       (.I0(\main_inst/main_float64_addexit_218_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_float64_addexit_218_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_float64_addexit_218_reg_reg_n_0_[14] ),
        .I3(\main_inst/main_float64_addexit_218_reg_reg_n_0_[15] ),
        .I4(\cur_state[1]_i_20_n_0 ),
        .O(\cur_state[1]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[1]_i_91 
       (.I0(\main_inst/main_15_19_reg [40]),
        .I1(\main_inst/main_15_19_reg [39]),
        .O(\cur_state[1]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_92 
       (.I0(\main_inst/main_15_19_reg [38]),
        .I1(\main_inst/main_15_19_reg [37]),
        .I2(\main_inst/main_15_19_reg [36]),
        .O(\cur_state[1]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_93 
       (.I0(\main_inst/main_15_19_reg [35]),
        .I1(\main_inst/main_15_19_reg [34]),
        .I2(\main_inst/main_15_19_reg [33]),
        .O(\cur_state[1]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_95 
       (.I0(\main_inst/main_15_19_reg [32]),
        .I1(\main_inst/main_15_19_reg [31]),
        .I2(\main_inst/main_15_19_reg [30]),
        .O(\cur_state[1]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_96 
       (.I0(\main_inst/main_15_19_reg [29]),
        .I1(\main_inst/main_15_19_reg [28]),
        .I2(\main_inst/main_15_19_reg [27]),
        .O(\cur_state[1]_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_97 
       (.I0(\main_inst/main_15_19_reg [26]),
        .I1(\main_inst/main_15_19_reg [25]),
        .I2(\main_inst/main_15_19_reg [24]),
        .O(\cur_state[1]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_98 
       (.I0(\main_inst/main_15_19_reg [23]),
        .I1(\main_inst/main_15_19_reg [22]),
        .I2(\main_inst/main_15_19_reg [21]),
        .O(\cur_state[1]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[1]_i_99 
       (.I0(\main_inst/main_15_19_reg [20]),
        .I1(\main_inst/main_15_19_reg [19]),
        .I2(\main_inst/main_15_19_reg [18]),
        .O(\cur_state[1]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \cur_state[1]_rep_i_1 
       (.I0(\cur_state[1]_i_2_n_0 ),
        .I1(\cur_state[1]_i_3_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\cur_state[1]_i_4_n_0 ),
        .I4(\cur_state[1]_i_5_n_0 ),
        .I5(\cur_state_reg[1]_i_6_n_0 ),
        .O(\cur_state[1]_rep_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30B833BB30B80088)) 
    \cur_state[2]_i_1 
       (.I0(\cur_state[2]_i_2_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\cur_state[2]_i_3_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\cur_state[2]_i_4_n_0 ),
        .O(\main_inst/next_state [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'h3C7C)) 
    \cur_state[2]_i_11 
       (.I0(\main_inst/main_112_114 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[2]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_16 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [30]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [31]),
        .O(\cur_state[2]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_19 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [28]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [29]),
        .O(\cur_state[2]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4FE0F0F0)) 
    \cur_state[2]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\cur_state[3]_i_5_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_20 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [26]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [27]),
        .O(\cur_state[2]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_21 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [24]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [25]),
        .O(\cur_state[2]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_22 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [22]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [23]),
        .O(\cur_state[2]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_24 
       (.I0(\main_inst/main_103_107_reg [41]),
        .I1(\main_inst/main_103_107_reg [40]),
        .I2(\main_inst/main_103_107_reg [39]),
        .O(\cur_state[2]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_25 
       (.I0(\main_inst/main_103_107_reg [38]),
        .I1(\main_inst/main_103_107_reg [37]),
        .I2(\main_inst/main_103_107_reg [36]),
        .O(\cur_state[2]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_26 
       (.I0(\main_inst/main_103_107_reg [35]),
        .I1(\main_inst/main_103_107_reg [34]),
        .I2(\main_inst/main_103_107_reg [33]),
        .O(\cur_state[2]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_28 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [20]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [21]),
        .O(\cur_state[2]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_29 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [18]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [19]),
        .O(\cur_state[2]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \cur_state[2]_i_3 
       (.I0(\cur_state[2]_i_5_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\cur_state[2]_i_6_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\cur_state[2]_i_7_n_0 ),
        .O(\cur_state[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_30 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [16]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [17]),
        .O(\cur_state[2]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_31 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [14]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [15]),
        .O(\cur_state[2]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_33 
       (.I0(\main_inst/main_103_107_reg [32]),
        .I1(\main_inst/main_103_107_reg [31]),
        .I2(\main_inst/main_103_107_reg [30]),
        .O(\cur_state[2]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_34 
       (.I0(\main_inst/main_103_107_reg [29]),
        .I1(\main_inst/main_103_107_reg [28]),
        .I2(\main_inst/main_103_107_reg [27]),
        .O(\cur_state[2]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_35 
       (.I0(\main_inst/main_103_107_reg [26]),
        .I1(\main_inst/main_103_107_reg [25]),
        .I2(\main_inst/main_103_107_reg [24]),
        .O(\cur_state[2]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_36 
       (.I0(\main_inst/main_103_107_reg [23]),
        .I1(\main_inst/main_103_107_reg [22]),
        .I2(\main_inst/main_103_107_reg [21]),
        .O(\cur_state[2]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_37 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [6]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [7]),
        .O(\cur_state[2]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_38 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [12]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [13]),
        .O(\cur_state[2]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_39 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [10]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [11]),
        .O(\cur_state[2]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA0CFAFCFAFCFAFC0)) 
    \cur_state[2]_i_4 
       (.I0(\cur_state[2]_i_8_n_0 ),
        .I1(\cur_state[2]_i_9_n_0 ),
        .I2(\cur_state[6]_i_11_n_0 ),
        .I3(\cur_state[6]_i_13_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_40 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [8]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [9]),
        .O(\cur_state[2]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \cur_state[2]_i_41 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [6]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [7]),
        .O(\cur_state[2]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_42 
       (.I0(\main_inst/main_103_107_reg [20]),
        .I1(\main_inst/main_103_107_reg [19]),
        .I2(\main_inst/main_103_107_reg [18]),
        .O(\cur_state[2]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_43 
       (.I0(\main_inst/main_103_107_reg [17]),
        .I1(\main_inst/main_103_107_reg [16]),
        .I2(\main_inst/main_103_107_reg [15]),
        .O(\cur_state[2]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[2]_i_44 
       (.I0(\main_inst/main_103_107_reg [14]),
        .I1(\main_inst/main_103_107_reg [13]),
        .I2(\main_inst/main_103_107_reg [12]),
        .O(\cur_state[2]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[2]_i_45 
       (.I0(\main_inst/main_103_107_reg [10]),
        .I1(\main_inst/main_103_107_reg [11]),
        .O(\cur_state[2]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h7C)) 
    \cur_state[2]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h76BB)) 
    \cur_state[2]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/main_127_128 ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7CCFFFFF7CCF0000)) 
    \cur_state[2]_i_7 
       (.I0(\main_inst/main_123_124 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\cur_state[2]_i_11_n_0 ),
        .O(\cur_state[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF0F50F030FF30)) 
    \cur_state[2]_i_8 
       (.I0(\main_inst/main_33_34 ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3CF2)) 
    \cur_state[2]_i_9 
       (.I0(\main_inst/main_81_83 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[2]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30B833BB30B80088)) 
    \cur_state[3]_i_1 
       (.I0(\cur_state[3]_i_2_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\cur_state_reg[3]_i_3_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\cur_state_reg[3]_i_4_n_0 ),
        .O(\main_inst/next_state [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hCCB0)) 
    \cur_state[3]_i_10 
       (.I0(\main_inst/main_112_114 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h5757AA8A)) 
    \cur_state[3]_i_13 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/main_23_24 ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\cur_state[3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h4C7CCCCC)) 
    \cur_state[3]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\cur_state[3]_i_5_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    \cur_state[3]_i_5 
       (.I0(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_4_n_0 ),
        .I1(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_5_n_0 ),
        .I2(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_6_n_0 ),
        .I3(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_7_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hDFFFFFFFDFFF0000)) 
    \cur_state[3]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/main_121_122 ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\cur_state[3]_i_10_n_0 ),
        .O(\cur_state[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h5FA0BABA)) 
    \cur_state[3]_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5DFFFFFF5DFF0000)) 
    \cur_state[3]_i_8 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2EAEEEAEEEAE2EAE)) 
    \cur_state[3]_i_9 
       (.I0(\cur_state[3]_i_13_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \cur_state[4]_i_1 
       (.I0(\cur_state[4]_i_2_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\cur_state[4]_i_3_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\cur_state[4]_i_4_n_0 ),
        .O(\main_inst/next_state [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4AAA0AAA0AAA0AAA)) 
    \cur_state[4]_i_2 
       (.I0(\cur_state[1]_i_5_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/main_float64_addexit_exitcond1_reg ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\cur_state[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB888)) 
    \cur_state[4]_i_3 
       (.I0(\cur_state[5]_i_4_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\cur_state[4]_i_5_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\cur_state[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFA0C0A0CFA0CFA0)) 
    \cur_state[4]_i_4 
       (.I0(\cur_state[4]_i_7_n_0 ),
        .I1(\cur_state[4]_i_8_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\cur_state[6]_i_12_n_0 ),
        .O(\cur_state[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \cur_state[4]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/main_123_124 ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \cur_state[4]_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0FC1)) 
    \cur_state[4]_i_8 
       (.I0(\main_inst/main_81_83 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[4]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000EEE22E22)) 
    \cur_state[5]_i_1 
       (.I0(\cur_state[5]_i_2_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\cur_state[5]_i_3_n_0 ),
        .I4(\cur_state[5]_i_4_n_0 ),
        .I5(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\cur_state[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_17 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .O(\cur_state[5]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_18 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .O(\cur_state[5]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_19 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .O(\cur_state[5]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000080)) 
    \cur_state[5]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_21 
       (.I0(\main_inst/main_103_107_reg [40]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_103_107_reg [41]),
        .O(\cur_state[5]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_22 
       (.I0(\main_inst/main_103_107_reg [38]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_103_107_reg [39]),
        .O(\cur_state[5]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_23 
       (.I0(\main_inst/main_103_107_reg [36]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_103_107_reg [37]),
        .O(\cur_state[5]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_24 
       (.I0(\main_inst/main_103_107_reg [34]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_103_107_reg [35]),
        .O(\cur_state[5]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_25 
       (.I0(\main_inst/main_103_107_reg [40]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_103_107_reg [41]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .O(\cur_state[5]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_26 
       (.I0(\main_inst/main_103_107_reg [38]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I2(\main_inst/main_103_107_reg [39]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .O(\cur_state[5]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_27 
       (.I0(\main_inst/main_103_107_reg [36]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_103_107_reg [37]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .O(\cur_state[5]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_28 
       (.I0(\main_inst/main_103_107_reg [34]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_103_107_reg [35]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .O(\cur_state[5]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFFFFFFF3FF00F0F)) 
    \cur_state[5]_i_3 
       (.I0(\main_inst/main_123_124 ),
        .I1(\main_inst/main_121_122 ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_30 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_103_107_reg [40]),
        .I2(\main_inst/main_103_107_reg [41]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .O(\cur_state[5]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_31 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_103_107_reg [38]),
        .I2(\main_inst/main_103_107_reg [39]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .O(\cur_state[5]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_32 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_103_107_reg [36]),
        .I2(\main_inst/main_103_107_reg [37]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .O(\cur_state[5]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_33 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_103_107_reg [34]),
        .I2(\main_inst/main_103_107_reg [35]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .O(\cur_state[5]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_34 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_103_107_reg [40]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_103_107_reg [41]),
        .O(\cur_state[5]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_35 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_103_107_reg [38]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_103_107_reg [39]),
        .O(\cur_state[5]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_36 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_103_107_reg [36]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_103_107_reg [37]),
        .O(\cur_state[5]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_37 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_103_107_reg [34]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_103_107_reg [35]),
        .O(\cur_state[5]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_39 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .O(\cur_state[5]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h3CFF334F)) 
    \cur_state[5]_i_4 
       (.I0(\main_inst/main_165_166 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_40 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .O(\cur_state[5]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_41 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .O(\cur_state[5]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_42 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .O(\cur_state[5]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_44 
       (.I0(\main_inst/main_103_107_reg [32]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_103_107_reg [33]),
        .O(\cur_state[5]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_45 
       (.I0(\main_inst/main_103_107_reg [30]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .I3(\main_inst/main_103_107_reg [31]),
        .O(\cur_state[5]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_46 
       (.I0(\main_inst/main_103_107_reg [28]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .I3(\main_inst/main_103_107_reg [29]),
        .O(\cur_state[5]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_47 
       (.I0(\main_inst/main_103_107_reg [26]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .I3(\main_inst/main_103_107_reg [27]),
        .O(\cur_state[5]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_48 
       (.I0(\main_inst/main_103_107_reg [32]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I2(\main_inst/main_103_107_reg [33]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .O(\cur_state[5]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_49 
       (.I0(\main_inst/main_103_107_reg [30]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I2(\main_inst/main_103_107_reg [31]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .O(\cur_state[5]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_50 
       (.I0(\main_inst/main_103_107_reg [28]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_103_107_reg [29]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .O(\cur_state[5]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_51 
       (.I0(\main_inst/main_103_107_reg [26]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_103_107_reg [27]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .O(\cur_state[5]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_53 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_103_107_reg [32]),
        .I2(\main_inst/main_103_107_reg [33]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .O(\cur_state[5]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_54 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_103_107_reg [30]),
        .I2(\main_inst/main_103_107_reg [31]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .O(\cur_state[5]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_55 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_103_107_reg [28]),
        .I2(\main_inst/main_103_107_reg [29]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .O(\cur_state[5]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_56 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_103_107_reg [26]),
        .I2(\main_inst/main_103_107_reg [27]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .O(\cur_state[5]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_57 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_103_107_reg [32]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_103_107_reg [33]),
        .O(\cur_state[5]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_58 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_103_107_reg [30]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .I3(\main_inst/main_103_107_reg [31]),
        .O(\cur_state[5]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_59 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_103_107_reg [28]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .I3(\main_inst/main_103_107_reg [29]),
        .O(\cur_state[5]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_60 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_103_107_reg [26]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .I3(\main_inst/main_103_107_reg [27]),
        .O(\cur_state[5]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_61 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .O(\cur_state[5]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_62 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .O(\cur_state[5]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \cur_state[5]_i_63 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .O(\cur_state[5]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \cur_state[5]_i_64 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .O(\cur_state[5]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_66 
       (.I0(\main_inst/main_103_107_reg [24]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .I3(\main_inst/main_103_107_reg [25]),
        .O(\cur_state[5]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_67 
       (.I0(\main_inst/main_103_107_reg [22]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_103_107_reg [23]),
        .O(\cur_state[5]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_68 
       (.I0(\main_inst/main_103_107_reg [20]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_103_107_reg [21]),
        .O(\cur_state[5]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_69 
       (.I0(\main_inst/main_103_107_reg [18]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_103_107_reg [19]),
        .O(\cur_state[5]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_70 
       (.I0(\main_inst/main_103_107_reg [24]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I2(\main_inst/main_103_107_reg [25]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .O(\cur_state[5]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_71 
       (.I0(\main_inst/main_103_107_reg [22]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_103_107_reg [23]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .O(\cur_state[5]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_72 
       (.I0(\main_inst/main_103_107_reg [20]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_103_107_reg [21]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .O(\cur_state[5]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_73 
       (.I0(\main_inst/main_103_107_reg [18]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I2(\main_inst/main_103_107_reg [19]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .O(\cur_state[5]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_75 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_103_107_reg [24]),
        .I2(\main_inst/main_103_107_reg [25]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .O(\cur_state[5]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_76 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I1(\main_inst/main_103_107_reg [22]),
        .I2(\main_inst/main_103_107_reg [23]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .O(\cur_state[5]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_77 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_103_107_reg [20]),
        .I2(\main_inst/main_103_107_reg [21]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .O(\cur_state[5]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_78 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I1(\main_inst/main_103_107_reg [18]),
        .I2(\main_inst/main_103_107_reg [19]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .O(\cur_state[5]_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_79 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_103_107_reg [24]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .I3(\main_inst/main_103_107_reg [25]),
        .O(\cur_state[5]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_80 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I1(\main_inst/main_103_107_reg [22]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_103_107_reg [23]),
        .O(\cur_state[5]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_81 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_103_107_reg [20]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_103_107_reg [21]),
        .O(\cur_state[5]_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_82 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I1(\main_inst/main_103_107_reg [18]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_103_107_reg [19]),
        .O(\cur_state[5]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_83 
       (.I0(\main_inst/main_103_107_reg [16]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_103_107_reg [17]),
        .O(\cur_state[5]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_84 
       (.I0(\main_inst/main_103_107_reg [14]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_103_107_reg [15]),
        .O(\cur_state[5]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_85 
       (.I0(\main_inst/main_103_107_reg [12]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_103_107_reg [13]),
        .O(\cur_state[5]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_86 
       (.I0(\main_inst/main_103_107_reg [10]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_103_107_reg [11]),
        .O(\cur_state[5]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_87 
       (.I0(\main_inst/main_103_107_reg [16]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_103_107_reg [17]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .O(\cur_state[5]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_88 
       (.I0(\main_inst/main_103_107_reg [14]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_103_107_reg [15]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .O(\cur_state[5]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_89 
       (.I0(\main_inst/main_103_107_reg [12]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I2(\main_inst/main_103_107_reg [13]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .O(\cur_state[5]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_90 
       (.I0(\main_inst/main_103_107_reg [10]),
        .I1(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I2(\main_inst/main_103_107_reg [11]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .O(\cur_state[5]_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_91 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_103_107_reg [16]),
        .I2(\main_inst/main_103_107_reg [17]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .O(\cur_state[5]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_92 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_103_107_reg [14]),
        .I2(\main_inst/main_103_107_reg [15]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .O(\cur_state[5]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_93 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_103_107_reg [12]),
        .I2(\main_inst/main_103_107_reg [13]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .O(\cur_state[5]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h2F02)) 
    \cur_state[5]_i_94 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I1(\main_inst/main_103_107_reg [10]),
        .I2(\main_inst/main_103_107_reg [11]),
        .I3(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .O(\cur_state[5]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_95 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_103_107_reg [16]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_103_107_reg [17]),
        .O(\cur_state[5]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_96 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_103_107_reg [14]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_103_107_reg [15]),
        .O(\cur_state[5]_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_97 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_103_107_reg [12]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_103_107_reg [13]),
        .O(\cur_state[5]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h9009)) 
    \cur_state[5]_i_98 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I1(\main_inst/main_103_107_reg [10]),
        .I2(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_103_107_reg [11]),
        .O(\cur_state[5]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00FF002E)) 
    \cur_state[6]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\cur_state[6]_i_3_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\cur_state[6]_i_4_n_0 ),
        .O(\main_inst/cur_state ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BB888888BB88B8)) 
    \cur_state[6]_i_10 
       (.I0(\cur_state[6]_i_16_n_0 ),
        .I1(\cur_state[6]_i_13_n_0 ),
        .I2(\main_inst/main_81_83 ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[6]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \cur_state[6]_i_11 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\cur_state[6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \cur_state[6]_i_12 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .O(\cur_state[6]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5D)) 
    \cur_state[6]_i_13 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\cur_state[6]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h50C000F0000F00F0)) 
    \cur_state[6]_i_14 
       (.I0(\main_inst/main_123_124 ),
        .I1(\main_inst/main_121_122 ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\cur_state[6]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hC3CC00B0)) 
    \cur_state[6]_i_15 
       (.I0(\main_inst/main_165_166 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[6]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00400022)) 
    \cur_state[6]_i_16 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/main_23_24 ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\cur_state[6]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    \cur_state[6]_i_21 
       (.I0(\main_inst/main_15_19_reg [40]),
        .I1(\main_inst/main_91_92 [40]),
        .I2(\main_inst/main_91_92 [39]),
        .I3(\main_inst/main_15_19_reg [39]),
        .O(\cur_state[6]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_22 
       (.I0(\main_inst/main_15_19_reg [38]),
        .I1(\main_inst/main_91_92 [38]),
        .I2(\main_inst/main_15_19_reg [37]),
        .I3(\main_inst/main_91_92 [37]),
        .I4(\main_inst/main_91_92 [36]),
        .I5(\main_inst/main_15_19_reg [36]),
        .O(\cur_state[6]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_23 
       (.I0(\main_inst/main_15_19_reg [35]),
        .I1(\main_inst/main_91_92 [35]),
        .I2(\main_inst/main_15_19_reg [34]),
        .I3(\main_inst/main_91_92 [34]),
        .I4(\main_inst/main_91_92 [33]),
        .I5(\main_inst/main_15_19_reg [33]),
        .O(\cur_state[6]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_25 
       (.I0(\main_inst/main_15_19_reg [32]),
        .I1(\main_inst/main_91_92 [32]),
        .I2(\main_inst/main_15_19_reg [31]),
        .I3(\main_inst/main_91_92 [31]),
        .I4(\main_inst/main_91_92 [30]),
        .I5(\main_inst/main_15_19_reg [30]),
        .O(\cur_state[6]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_26 
       (.I0(\main_inst/main_15_19_reg [29]),
        .I1(\main_inst/main_91_92 [29]),
        .I2(\main_inst/main_15_19_reg [28]),
        .I3(\main_inst/main_91_92 [28]),
        .I4(\main_inst/main_91_92 [27]),
        .I5(\main_inst/main_15_19_reg [27]),
        .O(\cur_state[6]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_27 
       (.I0(\main_inst/main_15_19_reg [26]),
        .I1(\main_inst/main_91_92 [26]),
        .I2(\main_inst/main_15_19_reg [25]),
        .I3(\main_inst/main_91_92 [25]),
        .I4(\main_inst/main_91_92 [24]),
        .I5(\main_inst/main_15_19_reg [24]),
        .O(\cur_state[6]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_28 
       (.I0(\main_inst/main_15_19_reg [23]),
        .I1(\main_inst/main_91_92 [23]),
        .I2(\main_inst/main_15_19_reg [22]),
        .I3(\main_inst/main_91_92 [22]),
        .I4(\main_inst/main_91_92 [21]),
        .I5(\main_inst/main_15_19_reg [21]),
        .O(\cur_state[6]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_29 
       (.I0(\main_inst/main_15_19_reg [20]),
        .I1(\main_inst/main_91_92 [20]),
        .I2(\main_inst/main_15_19_reg [19]),
        .I3(\main_inst/main_91_92 [19]),
        .I4(\main_inst/main_91_92 [18]),
        .I5(\main_inst/main_15_19_reg [18]),
        .O(\cur_state[6]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \cur_state[6]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\cur_state[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_30 
       (.I0(\main_inst/main_15_19_reg [17]),
        .I1(\main_inst/main_91_92 [17]),
        .I2(\main_inst/main_15_19_reg [16]),
        .I3(\main_inst/main_91_92 [16]),
        .I4(\main_inst/main_91_92 [15]),
        .I5(\main_inst/main_15_19_reg [15]),
        .O(\cur_state[6]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_31 
       (.I0(\main_inst/main_15_19_reg [14]),
        .I1(\main_inst/main_91_92 [14]),
        .I2(\main_inst/main_15_19_reg [13]),
        .I3(\main_inst/main_91_92 [13]),
        .I4(\main_inst/main_91_92 [12]),
        .I5(\main_inst/main_15_19_reg [12]),
        .O(\cur_state[6]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \cur_state[6]_i_32 
       (.I0(\main_inst/main_15_19_reg [11]),
        .I1(\main_inst/main_91_92 [11]),
        .I2(\main_inst/main_15_19_reg [10]),
        .I3(\main_inst/main_91_92 [10]),
        .I4(\main_inst/main_91_92 [9]),
        .I5(\main_inst/main_15_19_reg [9]),
        .O(\cur_state[6]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF454045404540)) 
    \cur_state[6]_i_4 
       (.I0(\cur_state[6]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_finish_reg_reg_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(start),
        .I4(\cur_state[6]_i_7_n_0 ),
        .I5(\cur_state[6]_i_8_n_0 ),
        .O(\cur_state[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888B888B8BBB888)) 
    \cur_state[6]_i_5 
       (.I0(\cur_state_reg[6]_i_9_n_0 ),
        .I1(\cur_state[1]_i_5_n_0 ),
        .I2(\cur_state[6]_i_10_n_0 ),
        .I3(\cur_state[6]_i_11_n_0 ),
        .I4(\cur_state[6]_i_12_n_0 ),
        .I5(\cur_state[6]_i_13_n_0 ),
        .O(\cur_state[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5F1FFFFF5F5FFFFF)) 
    \cur_state[6]_i_6 
       (.I0(\cur_state[1]_i_5_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/main_float64_addexit_exitcond1_reg ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\cur_state[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFB)) 
    \cur_state[6]_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_finish_reg_reg_n_0 ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\cur_state[6]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3333333337373736)) 
    \cur_state[6]_i_8 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\cur_state[6]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \cur_state_reg[0]_i_15 
       (.I0(\cur_state[0]_i_16_n_0 ),
        .I1(\cur_state[0]_i_17_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .O(cur_state_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF8 \cur_state_reg[0]_i_4 
       (.I0(\cur_state_reg[0]_i_7_n_0 ),
        .I1(\cur_state_reg[0]_i_8_n_0 ),
        .O(\cur_state_reg[0]_i_4_n_0 ),
        .S(\main_inst/cur_state_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[0]_i_5 
       (.I0(\cur_state[0]_i_9_n_0 ),
        .I1(cur_state),
        .O(\cur_state_reg[0]_i_5_n_0 ),
        .S(\cur_state[6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[0]_i_7 
       (.I0(\cur_state[0]_i_11_n_0 ),
        .I1(\cur_state[0]_i_12_n_0 ),
        .O(\cur_state_reg[0]_i_7_n_0 ),
        .S(\main_inst/cur_state_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[0]_i_8 
       (.I0(\cur_state[0]_i_13_n_0 ),
        .I1(\cur_state[0]_i_14_n_0 ),
        .O(\cur_state_reg[0]_i_8_n_0 ),
        .S(\main_inst/cur_state_reg_n_0_[3] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_11 
       (.CI(\cur_state_reg[1]_i_22_n_0 ),
        .CO({\cur_state_reg[1]_i_11_n_0 ,\cur_state_reg[1]_i_11_n_1 ,\cur_state_reg[1]_i_11_n_2 ,\main_inst/main_175_176 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_169_expDiff1ii_reg [31]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\cur_state[1]_i_23_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_22 
       (.CI(\cur_state_reg[1]_i_29_n_0 ),
        .CO({\cur_state_reg[1]_i_22_n_0 ,\cur_state_reg[1]_i_22_n_1 ,\cur_state_reg[1]_i_22_n_2 ,\cur_state_reg[1]_i_22_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_30_n_0 ,\cur_state[1]_i_31_n_0 ,\cur_state[1]_i_32_n_0 ,\cur_state[1]_i_33_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_24 
       (.CI(\cur_state_reg[1]_i_34_n_0 ),
        .CO({\cur_state_reg[1]_i_24_n_0 ,\cur_state_reg[1]_i_24_n_1 ,\main_inst/main_112_114 ,\cur_state_reg[1]_i_24_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \cur_state_reg[1]_i_26 
       (.I0(\cur_state[1]_i_41_n_0 ),
        .I1(\cur_state[1]_i_42_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\cur_state_reg[1]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_29 
       (.CI(\cur_state_reg[1]_i_43_n_0 ),
        .CO({\cur_state_reg[1]_i_29_n_0 ,\cur_state_reg[1]_i_29_n_1 ,\cur_state_reg[1]_i_29_n_2 ,\cur_state_reg[1]_i_29_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_44_n_0 ,\cur_state[1]_i_45_n_0 ,\cur_state[1]_i_46_n_0 ,\cur_state[1]_i_47_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_34 
       (.CI(\cur_state_reg[1]_i_48_n_0 ),
        .CO({\cur_state_reg[1]_i_34_n_0 ,\cur_state_reg[1]_i_34_n_1 ,\cur_state_reg[1]_i_34_n_2 ,\cur_state_reg[1]_i_34_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_43 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[1]_i_43_n_0 ,\cur_state_reg[1]_i_43_n_1 ,\cur_state_reg[1]_i_43_n_2 ,\cur_state_reg[1]_i_43_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\cur_state[1]_i_56_n_0 }),
        .S({\cur_state[1]_i_57_n_0 ,\cur_state[1]_i_58_n_0 ,\cur_state[1]_i_59_n_0 ,\cur_state[1]_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_48 
       (.CI(\cur_state_reg[1]_i_61_n_0 ),
        .CO({\cur_state_reg[1]_i_48_n_0 ,\cur_state_reg[1]_i_48_n_1 ,\cur_state_reg[1]_i_48_n_2 ,\cur_state_reg[1]_i_48_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\cur_state[1]_i_62_n_0 ,\cur_state[1]_i_63_n_0 ,\cur_state[1]_i_64_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_55 
       (.CI(\cur_state_reg[1]_i_72_n_0 ),
        .CO({\cur_state_reg[1]_i_55_n_0 ,\cur_state_reg[1]_i_55_n_1 ,\main_inst/data24 ,\cur_state_reg[1]_i_55_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[1]_i_6 
       (.I0(\cur_state[1]_i_16_n_0 ),
        .I1(\cur_state[1]_i_17_n_0 ),
        .O(\cur_state_reg[1]_i_6_n_0 ),
        .S(\cur_state[6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_61 
       (.CI(\cur_state_reg[1]_i_73_n_0 ),
        .CO({\cur_state_reg[1]_i_61_n_0 ,\cur_state_reg[1]_i_61_n_1 ,\cur_state_reg[1]_i_61_n_2 ,\cur_state_reg[1]_i_61_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_74_n_0 ,\cur_state[1]_i_75_n_0 ,\cur_state[1]_i_76_n_0 ,\cur_state[1]_i_77_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_72 
       (.CI(\cur_state_reg[1]_i_85_n_0 ),
        .CO({\cur_state_reg[1]_i_72_n_0 ,\cur_state_reg[1]_i_72_n_1 ,\cur_state_reg[1]_i_72_n_2 ,\cur_state_reg[1]_i_72_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_73 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[1]_i_73_n_0 ,\cur_state_reg[1]_i_73_n_1 ,\cur_state_reg[1]_i_73_n_2 ,\cur_state_reg[1]_i_73_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_86_n_0 ,\cur_state[1]_i_87_n_0 ,\cur_state[1]_i_88_n_0 ,\cur_state[1]_i_89_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_85 
       (.CI(\cur_state_reg[1]_i_90_n_0 ),
        .CO({\cur_state_reg[1]_i_85_n_0 ,\cur_state_reg[1]_i_85_n_1 ,\cur_state_reg[1]_i_85_n_2 ,\cur_state_reg[1]_i_85_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\cur_state[1]_i_91_n_0 ,\cur_state[1]_i_92_n_0 ,\cur_state[1]_i_93_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_90 
       (.CI(\cur_state_reg[1]_i_94_n_0 ),
        .CO({\cur_state_reg[1]_i_90_n_0 ,\cur_state_reg[1]_i_90_n_1 ,\cur_state_reg[1]_i_90_n_2 ,\cur_state_reg[1]_i_90_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_95_n_0 ,\cur_state[1]_i_96_n_0 ,\cur_state[1]_i_97_n_0 ,\cur_state[1]_i_98_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[1]_i_94 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[1]_i_94_n_0 ,\cur_state_reg[1]_i_94_n_1 ,\cur_state_reg[1]_i_94_n_2 ,\cur_state_reg[1]_i_94_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[1]_i_99_n_0 ,\cur_state[1]_i_100_n_0 ,\cur_state[1]_i_101_n_0 ,\cur_state[1]_i_102_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_10 
       (.CI(\cur_state_reg[2]_i_14_n_0 ),
        .CO({\cur_state_reg[2]_i_10_n_0 ,\cur_state_reg[2]_i_10_n_1 ,\main_inst/main_127_128 ,\cur_state_reg[2]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_12 
       (.CI(\cur_state_reg[2]_i_15_n_0 ),
        .CO({\cur_state_reg[2]_i_12_n_0 ,\cur_state_reg[2]_i_12_n_1 ,\cur_state_reg[2]_i_12_n_2 ,\main_inst/main_33_34 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_27_expDiff0i2i_reg [31]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\cur_state[2]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_14 
       (.CI(\cur_state_reg[2]_i_17_n_0 ),
        .CO({\cur_state_reg[2]_i_14_n_0 ,\cur_state_reg[2]_i_14_n_1 ,\cur_state_reg[2]_i_14_n_2 ,\cur_state_reg[2]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_15 
       (.CI(\cur_state_reg[2]_i_18_n_0 ),
        .CO({\cur_state_reg[2]_i_15_n_0 ,\cur_state_reg[2]_i_15_n_1 ,\cur_state_reg[2]_i_15_n_2 ,\cur_state_reg[2]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[2]_i_19_n_0 ,\cur_state[2]_i_20_n_0 ,\cur_state[2]_i_21_n_0 ,\cur_state[2]_i_22_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_17 
       (.CI(\cur_state_reg[2]_i_23_n_0 ),
        .CO({\cur_state_reg[2]_i_17_n_0 ,\cur_state_reg[2]_i_17_n_1 ,\cur_state_reg[2]_i_17_n_2 ,\cur_state_reg[2]_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\cur_state[2]_i_24_n_0 ,\cur_state[2]_i_25_n_0 ,\cur_state[2]_i_26_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_18 
       (.CI(\cur_state_reg[2]_i_27_n_0 ),
        .CO({\cur_state_reg[2]_i_18_n_0 ,\cur_state_reg[2]_i_18_n_1 ,\cur_state_reg[2]_i_18_n_2 ,\cur_state_reg[2]_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[2]_i_28_n_0 ,\cur_state[2]_i_29_n_0 ,\cur_state[2]_i_30_n_0 ,\cur_state[2]_i_31_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_23 
       (.CI(\cur_state_reg[2]_i_32_n_0 ),
        .CO({\cur_state_reg[2]_i_23_n_0 ,\cur_state_reg[2]_i_23_n_1 ,\cur_state_reg[2]_i_23_n_2 ,\cur_state_reg[2]_i_23_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[2]_i_33_n_0 ,\cur_state[2]_i_34_n_0 ,\cur_state[2]_i_35_n_0 ,\cur_state[2]_i_36_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_27 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[2]_i_27_n_0 ,\cur_state_reg[2]_i_27_n_1 ,\cur_state_reg[2]_i_27_n_2 ,\cur_state_reg[2]_i_27_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\cur_state[2]_i_37_n_0 }),
        .S({\cur_state[2]_i_38_n_0 ,\cur_state[2]_i_39_n_0 ,\cur_state[2]_i_40_n_0 ,\cur_state[2]_i_41_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[2]_i_32 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[2]_i_32_n_0 ,\cur_state_reg[2]_i_32_n_1 ,\cur_state_reg[2]_i_32_n_2 ,\cur_state_reg[2]_i_32_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[2]_i_42_n_0 ,\cur_state[2]_i_43_n_0 ,\cur_state[2]_i_44_n_0 ,\cur_state[2]_i_45_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[3]_i_3 
       (.I0(\cur_state[3]_i_6_n_0 ),
        .I1(\cur_state[3]_i_7_n_0 ),
        .O(\cur_state_reg[3]_i_3_n_0 ),
        .S(\main_inst/cur_state_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[3]_i_4 
       (.I0(\cur_state[3]_i_8_n_0 ),
        .I1(\cur_state[3]_i_9_n_0 ),
        .O(\cur_state_reg[3]_i_4_n_0 ),
        .S(\cur_state[6]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_10 
       (.CI(\cur_state_reg[5]_i_13_n_0 ),
        .CO({\cur_state_reg[5]_i_10_n_0 ,\cur_state_reg[5]_i_10_n_1 ,\cur_state_reg[5]_i_10_n_2 ,\cur_state_reg[5]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_11 
       (.CI(\cur_state_reg[5]_i_14_n_0 ),
        .CO({\cur_state_reg[5]_i_11_n_0 ,\cur_state_reg[5]_i_11_n_1 ,\cur_state_reg[5]_i_11_n_2 ,\cur_state_reg[5]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_12 
       (.CI(\cur_state_reg[5]_i_15_n_0 ),
        .CO({\cur_state_reg[5]_i_12_n_0 ,\cur_state_reg[5]_i_12_n_1 ,\cur_state_reg[5]_i_12_n_2 ,\cur_state_reg[5]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_13 
       (.CI(\cur_state_reg[5]_i_16_n_0 ),
        .CO({\cur_state_reg[5]_i_13_n_0 ,\cur_state_reg[5]_i_13_n_1 ,\cur_state_reg[5]_i_13_n_2 ,\cur_state_reg[5]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\cur_state[5]_i_17_n_0 ,\cur_state[5]_i_18_n_0 ,\cur_state[5]_i_19_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_14 
       (.CI(\cur_state_reg[5]_i_20_n_0 ),
        .CO({\cur_state_reg[5]_i_14_n_0 ,\cur_state_reg[5]_i_14_n_1 ,\cur_state_reg[5]_i_14_n_2 ,\cur_state_reg[5]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_21_n_0 ,\cur_state[5]_i_22_n_0 ,\cur_state[5]_i_23_n_0 ,\cur_state[5]_i_24_n_0 }),
        .S({\cur_state[5]_i_25_n_0 ,\cur_state[5]_i_26_n_0 ,\cur_state[5]_i_27_n_0 ,\cur_state[5]_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_15 
       (.CI(\cur_state_reg[5]_i_29_n_0 ),
        .CO({\cur_state_reg[5]_i_15_n_0 ,\cur_state_reg[5]_i_15_n_1 ,\cur_state_reg[5]_i_15_n_2 ,\cur_state_reg[5]_i_15_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_30_n_0 ,\cur_state[5]_i_31_n_0 ,\cur_state[5]_i_32_n_0 ,\cur_state[5]_i_33_n_0 }),
        .S({\cur_state[5]_i_34_n_0 ,\cur_state[5]_i_35_n_0 ,\cur_state[5]_i_36_n_0 ,\cur_state[5]_i_37_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_16 
       (.CI(\cur_state_reg[5]_i_38_n_0 ),
        .CO({\cur_state_reg[5]_i_16_n_0 ,\cur_state_reg[5]_i_16_n_1 ,\cur_state_reg[5]_i_16_n_2 ,\cur_state_reg[5]_i_16_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[5]_i_39_n_0 ,\cur_state[5]_i_40_n_0 ,\cur_state[5]_i_41_n_0 ,\cur_state[5]_i_42_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_20 
       (.CI(\cur_state_reg[5]_i_43_n_0 ),
        .CO({\cur_state_reg[5]_i_20_n_0 ,\cur_state_reg[5]_i_20_n_1 ,\cur_state_reg[5]_i_20_n_2 ,\cur_state_reg[5]_i_20_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_44_n_0 ,\cur_state[5]_i_45_n_0 ,\cur_state[5]_i_46_n_0 ,\cur_state[5]_i_47_n_0 }),
        .S({\cur_state[5]_i_48_n_0 ,\cur_state[5]_i_49_n_0 ,\cur_state[5]_i_50_n_0 ,\cur_state[5]_i_51_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_29 
       (.CI(\cur_state_reg[5]_i_52_n_0 ),
        .CO({\cur_state_reg[5]_i_29_n_0 ,\cur_state_reg[5]_i_29_n_1 ,\cur_state_reg[5]_i_29_n_2 ,\cur_state_reg[5]_i_29_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_53_n_0 ,\cur_state[5]_i_54_n_0 ,\cur_state[5]_i_55_n_0 ,\cur_state[5]_i_56_n_0 }),
        .S({\cur_state[5]_i_57_n_0 ,\cur_state[5]_i_58_n_0 ,\cur_state[5]_i_59_n_0 ,\cur_state[5]_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_38 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[5]_i_38_n_0 ,\cur_state_reg[5]_i_38_n_1 ,\cur_state_reg[5]_i_38_n_2 ,\cur_state_reg[5]_i_38_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[5]_i_61_n_0 ,\cur_state[5]_i_62_n_0 ,\cur_state[5]_i_63_n_0 ,\cur_state[5]_i_64_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_43 
       (.CI(\cur_state_reg[5]_i_65_n_0 ),
        .CO({\cur_state_reg[5]_i_43_n_0 ,\cur_state_reg[5]_i_43_n_1 ,\cur_state_reg[5]_i_43_n_2 ,\cur_state_reg[5]_i_43_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_66_n_0 ,\cur_state[5]_i_67_n_0 ,\cur_state[5]_i_68_n_0 ,\cur_state[5]_i_69_n_0 }),
        .S({\cur_state[5]_i_70_n_0 ,\cur_state[5]_i_71_n_0 ,\cur_state[5]_i_72_n_0 ,\cur_state[5]_i_73_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_5 
       (.CI(\cur_state_reg[5]_i_8_n_0 ),
        .CO({\cur_state_reg[5]_i_5_n_0 ,\cur_state_reg[5]_i_5_n_1 ,\main_inst/main_123_124 ,\cur_state_reg[5]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_52 
       (.CI(\cur_state_reg[5]_i_74_n_0 ),
        .CO({\cur_state_reg[5]_i_52_n_0 ,\cur_state_reg[5]_i_52_n_1 ,\cur_state_reg[5]_i_52_n_2 ,\cur_state_reg[5]_i_52_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_75_n_0 ,\cur_state[5]_i_76_n_0 ,\cur_state[5]_i_77_n_0 ,\cur_state[5]_i_78_n_0 }),
        .S({\cur_state[5]_i_79_n_0 ,\cur_state[5]_i_80_n_0 ,\cur_state[5]_i_81_n_0 ,\cur_state[5]_i_82_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_6 
       (.CI(\cur_state_reg[5]_i_9_n_0 ),
        .CO({\cur_state_reg[5]_i_6_n_0 ,\cur_state_reg[5]_i_6_n_1 ,\main_inst/main_121_122 ,\cur_state_reg[5]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_65 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[5]_i_65_n_0 ,\cur_state_reg[5]_i_65_n_1 ,\cur_state_reg[5]_i_65_n_2 ,\cur_state_reg[5]_i_65_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_83_n_0 ,\cur_state[5]_i_84_n_0 ,\cur_state[5]_i_85_n_0 ,\cur_state[5]_i_86_n_0 }),
        .S({\cur_state[5]_i_87_n_0 ,\cur_state[5]_i_88_n_0 ,\cur_state[5]_i_89_n_0 ,\cur_state[5]_i_90_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_7 
       (.CI(\cur_state_reg[5]_i_10_n_0 ),
        .CO({\cur_state_reg[5]_i_7_n_0 ,\cur_state_reg[5]_i_7_n_1 ,\main_inst/main_165_166 ,\cur_state_reg[5]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_74 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[5]_i_74_n_0 ,\cur_state_reg[5]_i_74_n_1 ,\cur_state_reg[5]_i_74_n_2 ,\cur_state_reg[5]_i_74_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\cur_state[5]_i_91_n_0 ,\cur_state[5]_i_92_n_0 ,\cur_state[5]_i_93_n_0 ,\cur_state[5]_i_94_n_0 }),
        .S({\cur_state[5]_i_95_n_0 ,\cur_state[5]_i_96_n_0 ,\cur_state[5]_i_97_n_0 ,\cur_state[5]_i_98_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_8 
       (.CI(\cur_state_reg[5]_i_11_n_0 ),
        .CO({\cur_state_reg[5]_i_8_n_0 ,\cur_state_reg[5]_i_8_n_1 ,\cur_state_reg[5]_i_8_n_2 ,\cur_state_reg[5]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[5]_i_9 
       (.CI(\cur_state_reg[5]_i_12_n_0 ),
        .CO({\cur_state_reg[5]_i_9_n_0 ,\cur_state_reg[5]_i_9_n_1 ,\cur_state_reg[5]_i_9_n_2 ,\cur_state_reg[5]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[6]_i_17 
       (.CI(\cur_state_reg[6]_i_18_n_0 ),
        .CO({\cur_state_reg[6]_i_17_n_0 ,\cur_state_reg[6]_i_17_n_1 ,\main_inst/main_81_83 ,\cur_state_reg[6]_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[6]_i_18 
       (.CI(\cur_state_reg[6]_i_19_n_0 ),
        .CO({\cur_state_reg[6]_i_18_n_0 ,\cur_state_reg[6]_i_18_n_1 ,\cur_state_reg[6]_i_18_n_2 ,\cur_state_reg[6]_i_18_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[6]_i_19 
       (.CI(\cur_state_reg[6]_i_20_n_0 ),
        .CO({\cur_state_reg[6]_i_19_n_0 ,\cur_state_reg[6]_i_19_n_1 ,\cur_state_reg[6]_i_19_n_2 ,\cur_state_reg[6]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\cur_state[6]_i_21_n_0 ,\cur_state[6]_i_22_n_0 ,\cur_state[6]_i_23_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[6]_i_2 
       (.I0(\cur_state[6]_i_5_n_0 ),
        .I1(\cur_state[6]_i_6_n_0 ),
        .O(\main_inst/next_state [6]),
        .S(\main_inst/cur_state_reg_n_0_[6] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[6]_i_20 
       (.CI(\cur_state_reg[6]_i_24_n_0 ),
        .CO({\cur_state_reg[6]_i_20_n_0 ,\cur_state_reg[6]_i_20_n_1 ,\cur_state_reg[6]_i_20_n_2 ,\cur_state_reg[6]_i_20_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[6]_i_25_n_0 ,\cur_state[6]_i_26_n_0 ,\cur_state[6]_i_27_n_0 ,\cur_state[6]_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \cur_state_reg[6]_i_24 
       (.CI(\<const0>__0__0 ),
        .CO({\cur_state_reg[6]_i_24_n_0 ,\cur_state_reg[6]_i_24_n_1 ,\cur_state_reg[6]_i_24_n_2 ,\cur_state_reg[6]_i_24_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\cur_state[6]_i_29_n_0 ,\cur_state[6]_i_30_n_0 ,\cur_state[6]_i_31_n_0 ,\cur_state[6]_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  MUXF7 \cur_state_reg[6]_i_9 
       (.I0(\cur_state[6]_i_14_n_0 ),
        .I1(\cur_state[6]_i_15_n_0 ),
        .O(\cur_state_reg[6]_i_9_n_0 ),
        .S(\main_inst/cur_state_reg_n_0_[4] ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h0E)) 
    finish_i_1
       (.I0(finish),
        .I1(\return_val[31]_i_2_n_0 ),
        .I2(\return_val[31]_i_1_n_0 ),
        .O(finish_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \main_101_102_reg[63]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(main_103_105_reg),
        .O(\main_inst/main_101_102_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[11]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(main_101_zExp1ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[11]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[11]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[11]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[15]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[15]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[15]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[15]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[19]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[19]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[19]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[19]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[23]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[23]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[23]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[23]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[27]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[27]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[27]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[27]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80004000)) 
    \main_101_zExp1ii_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_101_zExp1ii_reg[31]_i_3_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_inst/main_101_zSig0i12i_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \main_101_zExp1ii_reg[31]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_101_zExp1ii_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[31]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[31]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[31]_i_6 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[31]_i_7 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[3]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[3]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[3]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[3]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[7]_i_2 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[7]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[7]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zExp1ii_reg[7]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zExp1ii_reg[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[11]_i_1 
       (.CI(\main_101_zExp1ii_reg_reg[7]_i_1_n_0 ),
        .CO(main_101_zExp1ii_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[11]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[11]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[11]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[11]_i_1_n_7 }),
        .S({main_101_zExp1ii_reg,\main_101_zExp1ii_reg[11]_i_3_n_0 ,\main_101_zExp1ii_reg[11]_i_4_n_0 ,\main_101_zExp1ii_reg[11]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[15]_i_1 
       (.CI(main_101_zExp1ii_reg_reg[3]),
        .CO({\main_101_zExp1ii_reg_reg[15]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[15]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[15]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[15]_i_2_n_0 ,\main_101_zExp1ii_reg[15]_i_3_n_0 ,\main_101_zExp1ii_reg[15]_i_4_n_0 ,\main_101_zExp1ii_reg[15]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[19]_i_1 
       (.CI(\main_101_zExp1ii_reg_reg[15]_i_1_n_0 ),
        .CO({\main_101_zExp1ii_reg_reg[19]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[19]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[19]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[19]_i_2_n_0 ,\main_101_zExp1ii_reg[19]_i_3_n_0 ,\main_101_zExp1ii_reg[19]_i_4_n_0 ,\main_101_zExp1ii_reg[19]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[23]_i_1 
       (.CI(\main_101_zExp1ii_reg_reg[19]_i_1_n_0 ),
        .CO({\main_101_zExp1ii_reg_reg[23]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[23]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[23]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[23]_i_2_n_0 ,\main_101_zExp1ii_reg[23]_i_3_n_0 ,\main_101_zExp1ii_reg[23]_i_4_n_0 ,\main_101_zExp1ii_reg[23]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[27]_i_1 
       (.CI(\main_101_zExp1ii_reg_reg[23]_i_1_n_0 ),
        .CO({\main_101_zExp1ii_reg_reg[27]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[27]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[27]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[27]_i_2_n_0 ,\main_101_zExp1ii_reg[27]_i_3_n_0 ,\main_101_zExp1ii_reg[27]_i_4_n_0 ,\main_101_zExp1ii_reg[27]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[31]_i_2 
       (.CI(\main_101_zExp1ii_reg_reg[27]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[31]_i_2_n_4 ,\main_101_zExp1ii_reg_reg[31]_i_2_n_5 ,\main_101_zExp1ii_reg_reg[31]_i_2_n_6 ,\main_101_zExp1ii_reg_reg[31]_i_2_n_7 }),
        .S({\main_101_zExp1ii_reg[31]_i_4_n_0 ,\main_101_zExp1ii_reg[31]_i_5_n_0 ,\main_101_zExp1ii_reg[31]_i_6_n_0 ,\main_101_zExp1ii_reg[31]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\main_101_zExp1ii_reg_reg[3]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[3]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[3]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[3]_i_2_n_0 ,\main_101_zExp1ii_reg[3]_i_3_n_0 ,\main_101_zExp1ii_reg[3]_i_4_n_0 ,\main_101_zExp1ii_reg[3]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zExp1ii_reg_reg[7]_i_1 
       (.CI(\main_101_zExp1ii_reg_reg[3]_i_1_n_0 ),
        .CO({\main_101_zExp1ii_reg_reg[7]_i_1_n_0 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_1 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_2 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zExp1ii_reg_reg[7]_i_1_n_4 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_5 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_6 ,\main_101_zExp1ii_reg_reg[7]_i_1_n_7 }),
        .S({\main_101_zExp1ii_reg[7]_i_2_n_0 ,\main_101_zExp1ii_reg[7]_i_3_n_0 ,\main_101_zExp1ii_reg[7]_i_4_n_0 ,\main_101_zExp1ii_reg[7]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[12]_i_2 
       (.I0(\main_inst/main_15_19_reg [12]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(main_101_zSig0i12i_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[12]_i_3 
       (.I0(\main_inst/main_15_19_reg [11]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[12]_i_4 
       (.I0(\main_inst/main_15_19_reg [10]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[12]_i_5 
       (.I0(\main_inst/main_15_19_reg [9]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[12]_i_6 
       (.I0(\main_inst/main_15_19_reg [12]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [12]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [12]),
        .O(\main_101_zSig0i12i_reg[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[12]_i_7 
       (.I0(\main_inst/main_15_19_reg [11]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [11]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [11]),
        .O(\main_101_zSig0i12i_reg[12]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[12]_i_8 
       (.I0(\main_inst/main_15_19_reg [10]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [10]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [10]),
        .O(\main_101_zSig0i12i_reg[12]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[12]_i_9 
       (.I0(\main_inst/main_15_19_reg [9]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [9]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [9]),
        .O(\main_101_zSig0i12i_reg[12]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[16]_i_2 
       (.I0(\main_inst/main_15_19_reg [16]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[16]_i_3 
       (.I0(\main_inst/main_15_19_reg [15]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[16]_i_4 
       (.I0(\main_inst/main_15_19_reg [14]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[16]_i_5 
       (.I0(\main_inst/main_15_19_reg [13]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[16]_i_6 
       (.I0(\main_inst/main_15_19_reg [16]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [16]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [16]),
        .O(\main_101_zSig0i12i_reg[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[16]_i_7 
       (.I0(\main_inst/main_15_19_reg [15]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [15]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [15]),
        .O(\main_101_zSig0i12i_reg[16]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[16]_i_8 
       (.I0(\main_inst/main_15_19_reg [14]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [14]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [14]),
        .O(\main_101_zSig0i12i_reg[16]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[16]_i_9 
       (.I0(\main_inst/main_15_19_reg [13]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [13]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [13]),
        .O(\main_101_zSig0i12i_reg[16]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[20]_i_2 
       (.I0(\main_inst/main_15_19_reg [20]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[20]_i_3 
       (.I0(\main_inst/main_15_19_reg [19]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[20]_i_4 
       (.I0(\main_inst/main_15_19_reg [18]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[20]_i_5 
       (.I0(\main_inst/main_15_19_reg [17]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[20]_i_6 
       (.I0(\main_inst/main_15_19_reg [20]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [20]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [20]),
        .O(\main_101_zSig0i12i_reg[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[20]_i_7 
       (.I0(\main_inst/main_15_19_reg [19]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [19]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [19]),
        .O(\main_101_zSig0i12i_reg[20]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[20]_i_8 
       (.I0(\main_inst/main_15_19_reg [18]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [18]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [18]),
        .O(\main_101_zSig0i12i_reg[20]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[20]_i_9 
       (.I0(\main_inst/main_15_19_reg [17]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [17]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [17]),
        .O(\main_101_zSig0i12i_reg[20]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[24]_i_2 
       (.I0(\main_inst/main_15_19_reg [24]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[24]_i_3 
       (.I0(\main_inst/main_15_19_reg [23]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[24]_i_4 
       (.I0(\main_inst/main_15_19_reg [22]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[24]_i_5 
       (.I0(\main_inst/main_15_19_reg [21]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[24]_i_6 
       (.I0(\main_inst/main_15_19_reg [24]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [24]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [24]),
        .O(\main_101_zSig0i12i_reg[24]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[24]_i_7 
       (.I0(\main_inst/main_15_19_reg [23]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [23]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [23]),
        .O(\main_101_zSig0i12i_reg[24]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[24]_i_8 
       (.I0(\main_inst/main_15_19_reg [22]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [22]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [22]),
        .O(\main_101_zSig0i12i_reg[24]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[24]_i_9 
       (.I0(\main_inst/main_15_19_reg [21]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [21]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [21]),
        .O(\main_101_zSig0i12i_reg[24]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[28]_i_2 
       (.I0(\main_inst/main_15_19_reg [28]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[28]_i_3 
       (.I0(\main_inst/main_15_19_reg [27]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[28]_i_4 
       (.I0(\main_inst/main_15_19_reg [26]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[28]_i_5 
       (.I0(\main_inst/main_15_19_reg [25]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[28]_i_6 
       (.I0(\main_inst/main_15_19_reg [28]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [28]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [28]),
        .O(\main_101_zSig0i12i_reg[28]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[28]_i_7 
       (.I0(\main_inst/main_15_19_reg [27]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [27]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [27]),
        .O(\main_101_zSig0i12i_reg[28]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[28]_i_8 
       (.I0(\main_inst/main_15_19_reg [26]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [26]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [26]),
        .O(\main_101_zSig0i12i_reg[28]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[28]_i_9 
       (.I0(\main_inst/main_15_19_reg [25]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [25]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [25]),
        .O(\main_101_zSig0i12i_reg[28]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[32]_i_2 
       (.I0(\main_inst/main_15_19_reg [32]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[32]_i_3 
       (.I0(\main_inst/main_15_19_reg [31]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[32]_i_4 
       (.I0(\main_inst/main_15_19_reg [30]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[32]_i_5 
       (.I0(\main_inst/main_15_19_reg [29]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[32]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[32]_i_6 
       (.I0(\main_inst/main_15_19_reg [32]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [32]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [32]),
        .O(\main_101_zSig0i12i_reg[32]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[32]_i_7 
       (.I0(\main_inst/main_15_19_reg [31]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [31]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [31]),
        .O(\main_101_zSig0i12i_reg[32]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[32]_i_8 
       (.I0(\main_inst/main_15_19_reg [30]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [30]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [30]),
        .O(\main_101_zSig0i12i_reg[32]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[32]_i_9 
       (.I0(\main_inst/main_15_19_reg [29]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [29]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [29]),
        .O(\main_101_zSig0i12i_reg[32]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[36]_i_2 
       (.I0(\main_inst/main_15_19_reg [36]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[36]_i_3 
       (.I0(\main_inst/main_15_19_reg [35]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[36]_i_4 
       (.I0(\main_inst/main_15_19_reg [34]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[36]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[36]_i_5 
       (.I0(\main_inst/main_15_19_reg [33]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[36]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[36]_i_6 
       (.I0(\main_inst/main_15_19_reg [36]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [36]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [36]),
        .O(\main_101_zSig0i12i_reg[36]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[36]_i_7 
       (.I0(\main_inst/main_15_19_reg [35]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [35]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [35]),
        .O(\main_101_zSig0i12i_reg[36]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[36]_i_8 
       (.I0(\main_inst/main_15_19_reg [34]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [34]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [34]),
        .O(\main_101_zSig0i12i_reg[36]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[36]_i_9 
       (.I0(\main_inst/main_15_19_reg [33]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [33]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [33]),
        .O(\main_101_zSig0i12i_reg[36]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[40]_i_2 
       (.I0(\main_inst/main_15_19_reg [40]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[40]_i_3 
       (.I0(\main_inst/main_15_19_reg [39]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[40]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[40]_i_4 
       (.I0(\main_inst/main_15_19_reg [38]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[40]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_101_zSig0i12i_reg[40]_i_5 
       (.I0(\main_inst/main_15_19_reg [37]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[40]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[40]_i_6 
       (.I0(\main_inst/main_15_19_reg [40]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [40]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [40]),
        .O(\main_101_zSig0i12i_reg[40]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[40]_i_7 
       (.I0(\main_inst/main_15_19_reg [39]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [39]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [39]),
        .O(\main_101_zSig0i12i_reg[40]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[40]_i_8 
       (.I0(\main_inst/main_15_19_reg [38]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [38]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [38]),
        .O(\main_101_zSig0i12i_reg[40]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[40]_i_9 
       (.I0(\main_inst/main_15_19_reg [37]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [37]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [37]),
        .O(\main_101_zSig0i12i_reg[40]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zSig0i12i_reg[44]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_ii_reg [43]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[44]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zSig0i12i_reg[44]_i_4 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_ii_reg [42]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[44]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_101_zSig0i12i_reg[44]_i_5 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_ii_reg [41]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[44]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \main_101_zSig0i12i_reg[63]_i_3 
       (.I0(\main_inst/main_shift64RightJammingexit9ii_ii_reg [62]),
        .I1(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[63]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8000400000000000)) 
    \main_101_zSig0i12i_reg[8]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_101_zExp1ii_reg[31]_i_3_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_inst/main_101_zExp1ii1 ),
        .O(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5CAC)) 
    \main_101_zSig0i12i_reg[9]_i_1 
       (.I0(\main_inst/main_15_19_reg [9]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_ii_reg [9]),
        .I2(\main_inst/main_101_zExp1ii1 ),
        .I3(\main_inst/main_91_92 [9]),
        .O(\main_101_zSig0i12i_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000040)) 
    \main_101_zSig0i12i_reg[9]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(main_158_160_reg),
        .O(\main_inst/main_101_zExp1ii1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[12]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(main_101_zSig0i12i_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({main_101_zSig0i12i_reg,\main_101_zSig0i12i_reg[12]_i_3_n_0 ,\main_101_zSig0i12i_reg[12]_i_4_n_0 ,\main_101_zSig0i12i_reg[12]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[12]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[12]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[12]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[12]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[12]_i_6_n_0 ,\main_101_zSig0i12i_reg[12]_i_7_n_0 ,\main_101_zSig0i12i_reg[12]_i_8_n_0 ,\main_101_zSig0i12i_reg[12]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[16]_i_1 
       (.CI(main_101_zSig0i12i_reg_reg[3]),
        .CO({\main_101_zSig0i12i_reg_reg[16]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[16]_i_2_n_0 ,\main_101_zSig0i12i_reg[16]_i_3_n_0 ,\main_101_zSig0i12i_reg[16]_i_4_n_0 ,\main_101_zSig0i12i_reg[16]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[16]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[16]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[16]_i_6_n_0 ,\main_101_zSig0i12i_reg[16]_i_7_n_0 ,\main_101_zSig0i12i_reg[16]_i_8_n_0 ,\main_101_zSig0i12i_reg[16]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[20]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[16]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[20]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[20]_i_2_n_0 ,\main_101_zSig0i12i_reg[20]_i_3_n_0 ,\main_101_zSig0i12i_reg[20]_i_4_n_0 ,\main_101_zSig0i12i_reg[20]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[20]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[20]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[20]_i_6_n_0 ,\main_101_zSig0i12i_reg[20]_i_7_n_0 ,\main_101_zSig0i12i_reg[20]_i_8_n_0 ,\main_101_zSig0i12i_reg[20]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[24]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[20]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[24]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[24]_i_2_n_0 ,\main_101_zSig0i12i_reg[24]_i_3_n_0 ,\main_101_zSig0i12i_reg[24]_i_4_n_0 ,\main_101_zSig0i12i_reg[24]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[24]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[24]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[24]_i_6_n_0 ,\main_101_zSig0i12i_reg[24]_i_7_n_0 ,\main_101_zSig0i12i_reg[24]_i_8_n_0 ,\main_101_zSig0i12i_reg[24]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[28]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[24]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[28]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[28]_i_2_n_0 ,\main_101_zSig0i12i_reg[28]_i_3_n_0 ,\main_101_zSig0i12i_reg[28]_i_4_n_0 ,\main_101_zSig0i12i_reg[28]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[28]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[28]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[28]_i_6_n_0 ,\main_101_zSig0i12i_reg[28]_i_7_n_0 ,\main_101_zSig0i12i_reg[28]_i_8_n_0 ,\main_101_zSig0i12i_reg[28]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[32]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[28]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[32]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[32]_i_2_n_0 ,\main_101_zSig0i12i_reg[32]_i_3_n_0 ,\main_101_zSig0i12i_reg[32]_i_4_n_0 ,\main_101_zSig0i12i_reg[32]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[32]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[32]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[32]_i_6_n_0 ,\main_101_zSig0i12i_reg[32]_i_7_n_0 ,\main_101_zSig0i12i_reg[32]_i_8_n_0 ,\main_101_zSig0i12i_reg[32]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[36]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[32]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[36]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[36]_i_2_n_0 ,\main_101_zSig0i12i_reg[36]_i_3_n_0 ,\main_101_zSig0i12i_reg[36]_i_4_n_0 ,\main_101_zSig0i12i_reg[36]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[36]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[36]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[36]_i_6_n_0 ,\main_101_zSig0i12i_reg[36]_i_7_n_0 ,\main_101_zSig0i12i_reg[36]_i_8_n_0 ,\main_101_zSig0i12i_reg[36]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[40]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[36]_i_1_n_0 ),
        .CO({\main_101_zSig0i12i_reg_reg[40]_i_1_n_0 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_1 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_2 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_101_zSig0i12i_reg[40]_i_2_n_0 ,\main_101_zSig0i12i_reg[40]_i_3_n_0 ,\main_101_zSig0i12i_reg[40]_i_4_n_0 ,\main_101_zSig0i12i_reg[40]_i_5_n_0 }),
        .O({\main_101_zSig0i12i_reg_reg[40]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[40]_i_1_n_7 }),
        .S({\main_101_zSig0i12i_reg[40]_i_6_n_0 ,\main_101_zSig0i12i_reg[40]_i_7_n_0 ,\main_101_zSig0i12i_reg[40]_i_8_n_0 ,\main_101_zSig0i12i_reg[40]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[44]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[40]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zSig0i12i_reg_reg[44]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[44]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[44]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[44]_i_1_n_7 }),
        .S({ZERO_234,\main_101_zSig0i12i_reg[44]_i_3_n_0 ,\main_101_zSig0i12i_reg[44]_i_4_n_0 ,\main_101_zSig0i12i_reg[44]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  GND \main_101_zSig0i12i_reg_reg[60]_i_1_GND 
       (.G(\main_101_zSig0i12i_reg_reg[60]_i_1_GND_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_101_zSig0i12i_reg_reg[63]_i_1 
       (.CI(\main_101_zSig0i12i_reg_reg[60]_i_1_GND_1 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_101_zSig0i12i_reg_reg[63]_i_1_n_4 ,\main_101_zSig0i12i_reg_reg[63]_i_1_n_5 ,\main_101_zSig0i12i_reg_reg[63]_i_1_n_6 ,\main_101_zSig0i12i_reg_reg[63]_i_1_n_7 }),
        .S({\<const0>__0__0 ,ZERO_228,\main_101_zSig0i12i_reg[63]_i_3_n_0 ,ZERO_227}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \main_103_105_reg[41]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(main_103_105_reg),
        .O(\main_inst/main_103_105_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \main_103_105_reg[41]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .O(main_103_105_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00400000)) 
    \main_121_aExp0ii_reg[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .I5(\main_inst/main_121_aExp0ii_reg ),
        .O(main_121_aExp0ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00400000)) 
    \main_121_bExp0ii_reg[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .I5(\main_inst/main_121_bExp0ii_reg_reg_n_0_ ),
        .O(main_121_bExp0ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000000000000000)) 
    \main_136_expDiff0ii_reg[31]_i_1 
       (.I0(main_136_expDiff0ii_reg),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_inst/main_136_139_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \main_136_expDiff0ii_reg[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .O(main_136_expDiff0ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_136_expDiff0ii_reg_reg[4]_i_1_VCC 
       (.P(main_136_expDiff0ii_reg_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[0]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [0]),
        .I1(\main_inst/main_158_160 ),
        .O(main_158_159_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[10]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_ ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [10]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[11]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [11]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[12]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [12]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[13]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [13]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[14]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [14]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[15]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [15]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[16]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [16]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[17]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [17]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[18]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [18]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[19]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [19]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair359" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[1]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [1]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[20]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [20]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[21]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [21]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[22]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [22]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[23]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [23]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[24]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [24]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[25]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [25]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[26]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [26]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[27]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [27]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[28]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [28]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair322" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[29]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [29]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair358" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[2]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [2]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair321" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[30]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [30]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair320" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[31]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [31]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair319" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[32]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [32]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair318" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[33]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [33]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair317" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[34]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [34]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair316" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[35]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [35]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair315" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[36]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [36]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair314" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[37]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [37]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair313" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[38]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [38]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair312" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[39]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [39]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[3]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [3]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair311" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[40]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [40]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair310" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_158_159_reg[41]_i_1 
       (.I0(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [41]),
        .I2(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_159 [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair360" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[4]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [4]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[5]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [5]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[6]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [6]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[7]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [7]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair372" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[8]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [8]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair371" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_158_159_reg[9]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [9]),
        .I1(\main_inst/main_158_160 ),
        .O(\main_158_159_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00400000FFFFFFFF)) 
    \main_158_160_reg[62]_i_1 
       (.I0(main_158_160_reg),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_158_160_reg[62]_i_4_n_0 ),
        .I5(\main_inst/main_158_160 ),
        .O(\main_inst/main_158_bExp1ii_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \main_158_160_reg[62]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .O(main_158_160_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_158_160_reg[62]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_158_160_reg[62]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF7FFFFFFFFFFFFFF)) 
    \main_158_160_reg[62]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/main_123_124 ),
        .O(\main_inst/main_158_160 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair370" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_158_bExp1ii_reg[0]_i_1 
       (.I0(\main_inst/main_158_160 ),
        .I1(\main_inst/main_121_bExp0ii_reg_reg_n_0_ ),
        .O(main_158_bExp1ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_15_19_reg[40]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\return_val[31]_i_4_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_inst/main_15_17_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0008000000000000)) 
    \main_169_expDiff1ii_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\return_val[31]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_inst/main_169_172_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[11]_i_1_VCC 
       (.P(main_169_expDiff1ii_reg_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[15]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[19]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[23]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[27]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[31]_i_2_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[3]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_169_expDiff1ii_reg_reg[7]_i_1_VCC 
       (.P(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h4F)) 
    \main_191_192_reg[62]_i_1 
       (.I0(main_191_192_reg),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_aExp1ii_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFBFFFF)) 
    \main_191_192_reg[62]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/cur_state_reg_n_0_[4] ),
        .O(main_191_192_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFF7FFFFFFFFFF)) 
    \main_191_192_reg[62]_i_4 
       (.I0(\main_inst/main_121_122 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_inst/main_191_192 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[0]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [0]),
        .I1(\main_inst/main_191_192 ),
        .O(main_191_193_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[10]_i_1 
       (.I0(\main_inst/main_103_107_reg [10]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [10]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[11]_i_1 
       (.I0(\main_inst/main_103_107_reg [11]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [11]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[12]_i_1 
       (.I0(\main_inst/main_103_107_reg [12]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [12]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[13]_i_1 
       (.I0(\main_inst/main_103_107_reg [13]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [13]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[14]_i_1 
       (.I0(\main_inst/main_103_107_reg [14]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [14]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[15]_i_1 
       (.I0(\main_inst/main_103_107_reg [15]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [15]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[16]_i_1 
       (.I0(\main_inst/main_103_107_reg [16]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [16]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[17]_i_1 
       (.I0(\main_inst/main_103_107_reg [17]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [17]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[18]_i_1 
       (.I0(\main_inst/main_103_107_reg [18]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [18]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[19]_i_1 
       (.I0(\main_inst/main_103_107_reg [19]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [19]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[1]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [1]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[20]_i_1 
       (.I0(\main_inst/main_103_107_reg [20]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [20]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[21]_i_1 
       (.I0(\main_inst/main_103_107_reg [21]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [21]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[22]_i_1 
       (.I0(\main_inst/main_103_107_reg [22]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [22]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[23]_i_1 
       (.I0(\main_inst/main_103_107_reg [23]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [23]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[24]_i_1 
       (.I0(\main_inst/main_103_107_reg [24]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [24]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[25]_i_1 
       (.I0(\main_inst/main_103_107_reg [25]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [25]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[26]_i_1 
       (.I0(\main_inst/main_103_107_reg [26]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [26]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[27]_i_1 
       (.I0(\main_inst/main_103_107_reg [27]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [27]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[28]_i_1 
       (.I0(\main_inst/main_103_107_reg [28]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [28]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[29]_i_1 
       (.I0(\main_inst/main_103_107_reg [29]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [29]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[2]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [2]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[30]_i_1 
       (.I0(\main_inst/main_103_107_reg [30]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [30]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[31]_i_1 
       (.I0(\main_inst/main_103_107_reg [31]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [31]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[32]_i_1 
       (.I0(\main_inst/main_103_107_reg [32]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [32]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[33]_i_1 
       (.I0(\main_inst/main_103_107_reg [33]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [33]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[34]_i_1 
       (.I0(\main_inst/main_103_107_reg [34]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [34]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[35]_i_1 
       (.I0(\main_inst/main_103_107_reg [35]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [35]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[36]_i_1 
       (.I0(\main_inst/main_103_107_reg [36]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [36]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[37]_i_1 
       (.I0(\main_inst/main_103_107_reg [37]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [37]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[38]_i_1 
       (.I0(\main_inst/main_103_107_reg [38]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [38]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[39]_i_1 
       (.I0(\main_inst/main_103_107_reg [39]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [39]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[3]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [3]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[40]_i_1 
       (.I0(\main_inst/main_103_107_reg [40]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [40]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_191_193_reg[41]_i_1 
       (.I0(\main_inst/main_103_107_reg [41]),
        .I1(\main_inst/main_shift64RightJammingexitii_z0iii_reg [41]),
        .I2(\main_inst/main_191_192 ),
        .O(\main_inst/main_191_193 [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[4]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [4]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[5]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [5]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair369" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[6]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [6]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair368" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[7]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [7]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair367" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[8]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [8]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair366" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_191_193_reg[9]_i_1 
       (.I0(\main_inst/main_shift64RightJammingexitii_z0iii_reg [9]),
        .I1(\main_inst/main_191_192 ),
        .O(\main_191_193_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair365" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_191_aExp1ii_reg[0]_i_1 
       (.I0(\main_inst/main_191_192 ),
        .I1(\main_inst/main_121_aExp0ii_reg ),
        .O(main_191_aExp1ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \main_195_0ii_reg[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_158_160_reg[62]_i_4_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(main_195_0ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_10
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[50] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[51] ),
        .O(main_195_197_reg_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_11
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[48] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[49] ),
        .O(main_195_197_reg_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_13
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ),
        .O(main_195_197_reg_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_14
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ),
        .O(main_195_197_reg_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_15
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ),
        .O(main_195_197_reg_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_16
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ),
        .O(main_195_197_reg_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_17
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ),
        .O(main_195_197_reg_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_18
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[39] ),
        .O(main_195_197_reg_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_19
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[37] ),
        .O(main_195_197_reg_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_20
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[35] ),
        .O(main_195_197_reg_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    main_195_197_reg_i_21
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ),
        .O(main_195_197_reg_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_3
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ),
        .O(main_195_197_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_4
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ),
        .O(main_195_197_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_5
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ),
        .O(main_195_197_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_6
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ),
        .O(main_195_197_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_8
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[54] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[55] ),
        .O(main_195_197_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    main_195_197_reg_i_9
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[52] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[53] ),
        .O(main_195_197_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 main_195_197_reg_reg_i_1
       (.CI(main_195_197_reg_reg_i_2_n_0),
        .CO({\main_inst/main_195_197 ,main_195_197_reg_reg_i_1_n_1,main_195_197_reg_reg_i_1_n_2,main_195_197_reg_reg_i_1_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({main_195_197_reg_i_3_n_0,main_195_197_reg_i_4_n_0,main_195_197_reg_i_5_n_0,main_195_197_reg_i_6_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 main_195_197_reg_reg_i_12
       (.CI(\<const0>__0__0 ),
        .CO({main_195_197_reg_reg_i_12_n_0,main_195_197_reg_reg_i_12_n_1,main_195_197_reg_reg_i_12_n_2,main_195_197_reg_reg_i_12_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,main_195_197_reg_i_17_n_0}),
        .S({main_195_197_reg_i_18_n_0,main_195_197_reg_i_19_n_0,main_195_197_reg_i_20_n_0,main_195_197_reg_i_21_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 main_195_197_reg_reg_i_2
       (.CI(main_195_197_reg_reg_i_7_n_0),
        .CO({main_195_197_reg_reg_i_2_n_0,main_195_197_reg_reg_i_2_n_1,main_195_197_reg_reg_i_2_n_2,main_195_197_reg_reg_i_2_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({main_195_197_reg_i_8_n_0,main_195_197_reg_i_9_n_0,main_195_197_reg_i_10_n_0,main_195_197_reg_i_11_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 main_195_197_reg_reg_i_7
       (.CI(main_195_197_reg_reg_i_12_n_0),
        .CO({main_195_197_reg_reg_i_7_n_0,main_195_197_reg_reg_i_7_n_1,main_195_197_reg_reg_i_7_n_2,main_195_197_reg_reg_i_7_n_3}),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({main_195_197_reg_i_13_n_0,main_195_197_reg_i_14_n_0,main_195_197_reg_i_15_n_0,main_195_197_reg_i_16_n_0}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    main_195_199_reg_i_1
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(main_103_105_reg),
        .O(\main_inst/main_195_196_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACFCA)) 
    main_195_199_reg_i_10
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[48] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[49] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .O(main_195_199_reg_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    main_195_199_reg_i_2
       (.I0(main_195_199_reg_i_3_n_0),
        .I1(main_195_199_reg_i_4_n_0),
        .I2(main_195_199_reg_i_5_n_0),
        .I3(main_195_199_reg_i_6_n_0),
        .O(\main_inst/main_195_199 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFAFFCACFFFFFFFF)) 
    main_195_199_reg_i_3
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ),
        .I5(main_195_199_reg_i_7_n_0),
        .O(main_195_199_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000500353)) 
    main_195_199_reg_i_4
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ),
        .I5(main_195_199_reg_i_8_n_0),
        .O(main_195_199_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000500353)) 
    main_195_199_reg_i_5
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[55] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[54] ),
        .I5(main_195_199_reg_i_9_n_0),
        .O(main_195_199_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000500353)) 
    main_195_199_reg_i_6
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[51] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[50] ),
        .I5(main_195_199_reg_i_10_n_0),
        .O(main_195_199_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053035)) 
    main_195_199_reg_i_7
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .O(main_195_199_reg_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACFCA)) 
    main_195_199_reg_i_8
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .O(main_195_199_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACFCA)) 
    main_195_199_reg_i_9
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[52] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_195_197 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[53] ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .O(main_195_199_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[24]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[25]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[26]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[27]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[28]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[29]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[30]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_200_reg[31]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_200 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[24]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[25]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[26]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[27]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[28]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[29]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[30]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_extracttiiii_reg[31]_i_1 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ),
        .I2(\main_inst/main_195_197 ),
        .O(\main_inst/main_195_asinkiiii [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFF00000200)) 
    \main_195_iiiii_reg[4]_i_1 
       (.I0(\main_inst/main_195_iiiii ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_195_iiiii_reg[4]_i_2_n_0 ),
        .I5(\main_inst/main_195_iiiii_reg ),
        .O(main_195_iiiii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hEFFF)) 
    \main_195_iiiii_reg[4]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_195_iiiii_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \main_195_zExp0ii_reg[0]_i_1 
       (.I0(\main_inst/main_158_bExp1ii_reg_reg_n_0_ ),
        .I1(\main_inst/main_191_aExp1ii_reg_reg_n_0_ ),
        .I2(main_195_0ii_reg),
        .O(\main_inst/main_195_zExp0ii ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_2 
       (.I0(\main_inst/main_158_159_reg [11]),
        .I1(\main_inst/main_191_193_reg [11]),
        .I2(main_195_0ii_reg),
        .O(main_195_zSig0ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_3 
       (.I0(\main_inst/main_158_159_reg [10]),
        .I1(\main_inst/main_191_193_reg [10]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_4 
       (.I0(\main_inst/main_158_159_reg [9]),
        .I1(\main_inst/main_191_193_reg [9]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_5 
       (.I0(\main_inst/main_158_159_reg [8]),
        .I1(\main_inst/main_191_193_reg [8]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[11]_i_6 
       (.I0(\main_inst/main_191_193_reg [11]),
        .I1(\main_inst/main_158_159_reg [11]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [11]),
        .I4(\main_inst/main_158_160_reg [11]),
        .O(\main_195_zSig0ii_reg[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[11]_i_7 
       (.I0(\main_inst/main_191_193_reg [10]),
        .I1(\main_inst/main_158_159_reg [10]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [10]),
        .I4(\main_inst/main_158_160_reg [10]),
        .O(\main_195_zSig0ii_reg[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_8 
       (.I0(\main_inst/main_158_159_reg [9]),
        .I1(\main_inst/main_191_193_reg [9]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[11]_i_9 
       (.I0(\main_inst/main_158_159_reg [8]),
        .I1(\main_inst/main_191_193_reg [8]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[15]_i_2 
       (.I0(\main_inst/main_158_159_reg [15]),
        .I1(\main_inst/main_191_193_reg [15]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[15]_i_3 
       (.I0(\main_inst/main_158_159_reg [14]),
        .I1(\main_inst/main_191_193_reg [14]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[15]_i_4 
       (.I0(\main_inst/main_158_159_reg [13]),
        .I1(\main_inst/main_191_193_reg [13]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[15]_i_5 
       (.I0(\main_inst/main_158_159_reg [12]),
        .I1(\main_inst/main_191_193_reg [12]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[15]_i_6 
       (.I0(\main_inst/main_191_193_reg [15]),
        .I1(\main_inst/main_158_159_reg [15]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [15]),
        .I4(\main_inst/main_158_160_reg [15]),
        .O(\main_195_zSig0ii_reg[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[15]_i_7 
       (.I0(\main_inst/main_191_193_reg [14]),
        .I1(\main_inst/main_158_159_reg [14]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [14]),
        .I4(\main_inst/main_158_160_reg [14]),
        .O(\main_195_zSig0ii_reg[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[15]_i_8 
       (.I0(\main_inst/main_191_193_reg [13]),
        .I1(\main_inst/main_158_159_reg [13]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [13]),
        .I4(\main_inst/main_158_160_reg [13]),
        .O(\main_195_zSig0ii_reg[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[15]_i_9 
       (.I0(\main_inst/main_191_193_reg [12]),
        .I1(\main_inst/main_158_159_reg [12]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [12]),
        .I4(\main_inst/main_158_160_reg [12]),
        .O(\main_195_zSig0ii_reg[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[19]_i_2 
       (.I0(\main_inst/main_158_159_reg [19]),
        .I1(\main_inst/main_191_193_reg [19]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[19]_i_3 
       (.I0(\main_inst/main_158_159_reg [18]),
        .I1(\main_inst/main_191_193_reg [18]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[19]_i_4 
       (.I0(\main_inst/main_158_159_reg [17]),
        .I1(\main_inst/main_191_193_reg [17]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[19]_i_5 
       (.I0(\main_inst/main_158_159_reg [16]),
        .I1(\main_inst/main_191_193_reg [16]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[19]_i_6 
       (.I0(\main_inst/main_191_193_reg [19]),
        .I1(\main_inst/main_158_159_reg [19]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [19]),
        .I4(\main_inst/main_158_160_reg [19]),
        .O(\main_195_zSig0ii_reg[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[19]_i_7 
       (.I0(\main_inst/main_191_193_reg [18]),
        .I1(\main_inst/main_158_159_reg [18]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [18]),
        .I4(\main_inst/main_158_160_reg [18]),
        .O(\main_195_zSig0ii_reg[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[19]_i_8 
       (.I0(\main_inst/main_191_193_reg [17]),
        .I1(\main_inst/main_158_159_reg [17]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [17]),
        .I4(\main_inst/main_158_160_reg [17]),
        .O(\main_195_zSig0ii_reg[19]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[19]_i_9 
       (.I0(\main_inst/main_191_193_reg [16]),
        .I1(\main_inst/main_158_159_reg [16]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [16]),
        .I4(\main_inst/main_158_160_reg [16]),
        .O(\main_195_zSig0ii_reg[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[23]_i_2 
       (.I0(\main_inst/main_158_159_reg [23]),
        .I1(\main_inst/main_191_193_reg [23]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[23]_i_3 
       (.I0(\main_inst/main_158_159_reg [22]),
        .I1(\main_inst/main_191_193_reg [22]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[23]_i_4 
       (.I0(\main_inst/main_158_159_reg [21]),
        .I1(\main_inst/main_191_193_reg [21]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[23]_i_5 
       (.I0(\main_inst/main_158_159_reg [20]),
        .I1(\main_inst/main_191_193_reg [20]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[23]_i_6 
       (.I0(\main_inst/main_191_193_reg [23]),
        .I1(\main_inst/main_158_159_reg [23]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [23]),
        .I4(\main_inst/main_158_160_reg [23]),
        .O(\main_195_zSig0ii_reg[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[23]_i_7 
       (.I0(\main_inst/main_191_193_reg [22]),
        .I1(\main_inst/main_158_159_reg [22]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [22]),
        .I4(\main_inst/main_158_160_reg [22]),
        .O(\main_195_zSig0ii_reg[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[23]_i_8 
       (.I0(\main_inst/main_191_193_reg [21]),
        .I1(\main_inst/main_158_159_reg [21]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [21]),
        .I4(\main_inst/main_158_160_reg [21]),
        .O(\main_195_zSig0ii_reg[23]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[23]_i_9 
       (.I0(\main_inst/main_191_193_reg [20]),
        .I1(\main_inst/main_158_159_reg [20]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [20]),
        .I4(\main_inst/main_158_160_reg [20]),
        .O(\main_195_zSig0ii_reg[23]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[27]_i_2 
       (.I0(\main_inst/main_158_159_reg [27]),
        .I1(\main_inst/main_191_193_reg [27]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[27]_i_3 
       (.I0(\main_inst/main_158_159_reg [26]),
        .I1(\main_inst/main_191_193_reg [26]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[27]_i_4 
       (.I0(\main_inst/main_158_159_reg [25]),
        .I1(\main_inst/main_191_193_reg [25]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[27]_i_5 
       (.I0(\main_inst/main_158_159_reg [24]),
        .I1(\main_inst/main_191_193_reg [24]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[27]_i_6 
       (.I0(\main_inst/main_191_193_reg [27]),
        .I1(\main_inst/main_158_159_reg [27]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [27]),
        .I4(\main_inst/main_158_160_reg [27]),
        .O(\main_195_zSig0ii_reg[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[27]_i_7 
       (.I0(\main_inst/main_191_193_reg [26]),
        .I1(\main_inst/main_158_159_reg [26]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [26]),
        .I4(\main_inst/main_158_160_reg [26]),
        .O(\main_195_zSig0ii_reg[27]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[27]_i_8 
       (.I0(\main_inst/main_191_193_reg [25]),
        .I1(\main_inst/main_158_159_reg [25]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [25]),
        .I4(\main_inst/main_158_160_reg [25]),
        .O(\main_195_zSig0ii_reg[27]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[27]_i_9 
       (.I0(\main_inst/main_191_193_reg [24]),
        .I1(\main_inst/main_158_159_reg [24]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [24]),
        .I4(\main_inst/main_158_160_reg [24]),
        .O(\main_195_zSig0ii_reg[27]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[31]_i_2 
       (.I0(\main_inst/main_158_159_reg [31]),
        .I1(\main_inst/main_191_193_reg [31]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[31]_i_3 
       (.I0(\main_inst/main_158_159_reg [30]),
        .I1(\main_inst/main_191_193_reg [30]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[31]_i_4 
       (.I0(\main_inst/main_158_159_reg [29]),
        .I1(\main_inst/main_191_193_reg [29]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[31]_i_5 
       (.I0(\main_inst/main_158_159_reg [28]),
        .I1(\main_inst/main_191_193_reg [28]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[31]_i_6 
       (.I0(\main_inst/main_191_193_reg [31]),
        .I1(\main_inst/main_158_159_reg [31]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [31]),
        .I4(\main_inst/main_158_160_reg [31]),
        .O(\main_195_zSig0ii_reg[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[31]_i_7 
       (.I0(\main_inst/main_191_193_reg [30]),
        .I1(\main_inst/main_158_159_reg [30]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [30]),
        .I4(\main_inst/main_158_160_reg [30]),
        .O(\main_195_zSig0ii_reg[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[31]_i_8 
       (.I0(\main_inst/main_191_193_reg [29]),
        .I1(\main_inst/main_158_159_reg [29]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [29]),
        .I4(\main_inst/main_158_160_reg [29]),
        .O(\main_195_zSig0ii_reg[31]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[31]_i_9 
       (.I0(\main_inst/main_191_193_reg [28]),
        .I1(\main_inst/main_158_159_reg [28]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [28]),
        .I4(\main_inst/main_158_160_reg [28]),
        .O(\main_195_zSig0ii_reg[31]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[35]_i_2 
       (.I0(\main_inst/main_158_159_reg [35]),
        .I1(\main_inst/main_191_193_reg [35]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[35]_i_3 
       (.I0(\main_inst/main_158_159_reg [34]),
        .I1(\main_inst/main_191_193_reg [34]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[35]_i_4 
       (.I0(\main_inst/main_158_159_reg [33]),
        .I1(\main_inst/main_191_193_reg [33]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[35]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[35]_i_5 
       (.I0(\main_inst/main_158_159_reg [32]),
        .I1(\main_inst/main_191_193_reg [32]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[35]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[35]_i_6 
       (.I0(\main_inst/main_191_193_reg [35]),
        .I1(\main_inst/main_158_159_reg [35]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [35]),
        .I4(\main_inst/main_158_160_reg [35]),
        .O(\main_195_zSig0ii_reg[35]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[35]_i_7 
       (.I0(\main_inst/main_191_193_reg [34]),
        .I1(\main_inst/main_158_159_reg [34]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [34]),
        .I4(\main_inst/main_158_160_reg [34]),
        .O(\main_195_zSig0ii_reg[35]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[35]_i_8 
       (.I0(\main_inst/main_191_193_reg [33]),
        .I1(\main_inst/main_158_159_reg [33]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [33]),
        .I4(\main_inst/main_158_160_reg [33]),
        .O(\main_195_zSig0ii_reg[35]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[35]_i_9 
       (.I0(\main_inst/main_191_193_reg [32]),
        .I1(\main_inst/main_158_159_reg [32]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [32]),
        .I4(\main_inst/main_158_160_reg [32]),
        .O(\main_195_zSig0ii_reg[35]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[39]_i_2 
       (.I0(\main_inst/main_158_159_reg [39]),
        .I1(\main_inst/main_191_193_reg [39]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[39]_i_3 
       (.I0(\main_inst/main_158_159_reg [38]),
        .I1(\main_inst/main_191_193_reg [38]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[39]_i_4 
       (.I0(\main_inst/main_158_159_reg [37]),
        .I1(\main_inst/main_191_193_reg [37]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[39]_i_5 
       (.I0(\main_inst/main_158_159_reg [36]),
        .I1(\main_inst/main_191_193_reg [36]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[39]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[39]_i_6 
       (.I0(\main_inst/main_191_193_reg [39]),
        .I1(\main_inst/main_158_159_reg [39]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [39]),
        .I4(\main_inst/main_158_160_reg [39]),
        .O(\main_195_zSig0ii_reg[39]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[39]_i_7 
       (.I0(\main_inst/main_191_193_reg [38]),
        .I1(\main_inst/main_158_159_reg [38]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [38]),
        .I4(\main_inst/main_158_160_reg [38]),
        .O(\main_195_zSig0ii_reg[39]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[39]_i_8 
       (.I0(\main_inst/main_191_193_reg [37]),
        .I1(\main_inst/main_158_159_reg [37]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [37]),
        .I4(\main_inst/main_158_160_reg [37]),
        .O(\main_195_zSig0ii_reg[39]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[39]_i_9 
       (.I0(\main_inst/main_191_193_reg [36]),
        .I1(\main_inst/main_158_159_reg [36]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [36]),
        .I4(\main_inst/main_158_160_reg [36]),
        .O(\main_195_zSig0ii_reg[39]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_2 
       (.I0(\main_inst/main_158_159_reg [3]),
        .I1(\main_inst/main_191_193_reg [3]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_3 
       (.I0(\main_inst/main_158_159_reg [2]),
        .I1(\main_inst/main_191_193_reg [2]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_4 
       (.I0(\main_inst/main_158_159_reg [1]),
        .I1(\main_inst/main_191_193_reg [1]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_5 
       (.I0(\main_inst/main_158_159_reg [0]),
        .I1(\main_inst/main_191_193_reg [0]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_6 
       (.I0(\main_inst/main_158_159_reg [3]),
        .I1(\main_inst/main_191_193_reg [3]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_7 
       (.I0(\main_inst/main_158_159_reg [2]),
        .I1(\main_inst/main_191_193_reg [2]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_8 
       (.I0(\main_inst/main_158_159_reg [1]),
        .I1(\main_inst/main_191_193_reg [1]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[3]_i_9 
       (.I0(\main_inst/main_158_159_reg [0]),
        .I1(\main_inst/main_191_193_reg [0]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[43]_i_2 
       (.I0(\main_inst/main_158_159_reg [41]),
        .I1(\main_inst/main_191_193_reg [41]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[43]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[43]_i_3 
       (.I0(\main_inst/main_158_159_reg [40]),
        .I1(\main_inst/main_191_193_reg [40]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[43]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[43]_i_4 
       (.I0(\main_inst/main_191_193_reg [41]),
        .I1(\main_inst/main_158_159_reg [41]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [41]),
        .I4(\main_inst/main_158_160_reg [41]),
        .O(\main_195_zSig0ii_reg[43]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCAC53A35)) 
    \main_195_zSig0ii_reg[43]_i_5 
       (.I0(\main_inst/main_191_193_reg [40]),
        .I1(\main_inst/main_158_159_reg [40]),
        .I2(main_195_0ii_reg),
        .I3(\main_inst/main_191_192_reg [40]),
        .I4(\main_inst/main_158_160_reg [40]),
        .O(\main_195_zSig0ii_reg[43]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hF1)) 
    \main_195_zSig0ii_reg[63]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_195_zSig0ii_reg[63]_i_3_n_0 ),
        .I2(main_195_0ii_reg),
        .O(\main_inst/main_195_zSig0ii_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEFFFFFFFFFF)) 
    \main_195_zSig0ii_reg[63]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_195_zSig0ii_reg[63]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1B)) 
    \main_195_zSig0ii_reg[63]_i_4 
       (.I0(main_195_0ii_reg),
        .I1(\main_inst/main_191_192_reg [62]),
        .I2(\main_inst/main_158_160_reg [62]),
        .O(\main_195_zSig0ii_reg[63]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_2 
       (.I0(\main_inst/main_158_159_reg [7]),
        .I1(\main_inst/main_191_193_reg [7]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_3 
       (.I0(\main_inst/main_158_159_reg [6]),
        .I1(\main_inst/main_191_193_reg [6]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_4 
       (.I0(\main_inst/main_158_159_reg [5]),
        .I1(\main_inst/main_191_193_reg [5]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_5 
       (.I0(\main_inst/main_158_159_reg [4]),
        .I1(\main_inst/main_191_193_reg [4]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_6 
       (.I0(\main_inst/main_158_159_reg [7]),
        .I1(\main_inst/main_191_193_reg [7]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_7 
       (.I0(\main_inst/main_158_159_reg [6]),
        .I1(\main_inst/main_191_193_reg [6]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_8 
       (.I0(\main_inst/main_158_159_reg [5]),
        .I1(\main_inst/main_191_193_reg [5]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h53)) 
    \main_195_zSig0ii_reg[7]_i_9 
       (.I0(\main_inst/main_158_159_reg [4]),
        .I1(\main_inst/main_191_193_reg [4]),
        .I2(main_195_0ii_reg),
        .O(\main_195_zSig0ii_reg[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[11]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[7]_i_1_n_0 ),
        .CO(main_195_zSig0ii_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({main_195_zSig0ii_reg,\main_195_zSig0ii_reg[11]_i_3_n_0 ,\main_195_zSig0ii_reg[11]_i_4_n_0 ,\main_195_zSig0ii_reg[11]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [11:8]),
        .S({\main_195_zSig0ii_reg[11]_i_6_n_0 ,\main_195_zSig0ii_reg[11]_i_7_n_0 ,\main_195_zSig0ii_reg[11]_i_8_n_0 ,\main_195_zSig0ii_reg[11]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[15]_i_1 
       (.CI(main_195_zSig0ii_reg_reg[3]),
        .CO({\main_195_zSig0ii_reg_reg[15]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[15]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[15]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[15]_i_2_n_0 ,\main_195_zSig0ii_reg[15]_i_3_n_0 ,\main_195_zSig0ii_reg[15]_i_4_n_0 ,\main_195_zSig0ii_reg[15]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [15:12]),
        .S({\main_195_zSig0ii_reg[15]_i_6_n_0 ,\main_195_zSig0ii_reg[15]_i_7_n_0 ,\main_195_zSig0ii_reg[15]_i_8_n_0 ,\main_195_zSig0ii_reg[15]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[19]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[15]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[19]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[19]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[19]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[19]_i_2_n_0 ,\main_195_zSig0ii_reg[19]_i_3_n_0 ,\main_195_zSig0ii_reg[19]_i_4_n_0 ,\main_195_zSig0ii_reg[19]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [19:16]),
        .S({\main_195_zSig0ii_reg[19]_i_6_n_0 ,\main_195_zSig0ii_reg[19]_i_7_n_0 ,\main_195_zSig0ii_reg[19]_i_8_n_0 ,\main_195_zSig0ii_reg[19]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[23]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[19]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[23]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[23]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[23]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[23]_i_2_n_0 ,\main_195_zSig0ii_reg[23]_i_3_n_0 ,\main_195_zSig0ii_reg[23]_i_4_n_0 ,\main_195_zSig0ii_reg[23]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [23:20]),
        .S({\main_195_zSig0ii_reg[23]_i_6_n_0 ,\main_195_zSig0ii_reg[23]_i_7_n_0 ,\main_195_zSig0ii_reg[23]_i_8_n_0 ,\main_195_zSig0ii_reg[23]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[27]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[23]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[27]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[27]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[27]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[27]_i_2_n_0 ,\main_195_zSig0ii_reg[27]_i_3_n_0 ,\main_195_zSig0ii_reg[27]_i_4_n_0 ,\main_195_zSig0ii_reg[27]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [27:24]),
        .S({\main_195_zSig0ii_reg[27]_i_6_n_0 ,\main_195_zSig0ii_reg[27]_i_7_n_0 ,\main_195_zSig0ii_reg[27]_i_8_n_0 ,\main_195_zSig0ii_reg[27]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[31]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[27]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[31]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[31]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[31]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[31]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[31]_i_2_n_0 ,\main_195_zSig0ii_reg[31]_i_3_n_0 ,\main_195_zSig0ii_reg[31]_i_4_n_0 ,\main_195_zSig0ii_reg[31]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [31:28]),
        .S({\main_195_zSig0ii_reg[31]_i_6_n_0 ,\main_195_zSig0ii_reg[31]_i_7_n_0 ,\main_195_zSig0ii_reg[31]_i_8_n_0 ,\main_195_zSig0ii_reg[31]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[35]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[31]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[35]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[35]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[35]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[35]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[35]_i_2_n_0 ,\main_195_zSig0ii_reg[35]_i_3_n_0 ,\main_195_zSig0ii_reg[35]_i_4_n_0 ,\main_195_zSig0ii_reg[35]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [35:32]),
        .S({\main_195_zSig0ii_reg[35]_i_6_n_0 ,\main_195_zSig0ii_reg[35]_i_7_n_0 ,\main_195_zSig0ii_reg[35]_i_8_n_0 ,\main_195_zSig0ii_reg[35]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[39]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[35]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[39]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[39]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[39]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[39]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[39]_i_2_n_0 ,\main_195_zSig0ii_reg[39]_i_3_n_0 ,\main_195_zSig0ii_reg[39]_i_4_n_0 ,\main_195_zSig0ii_reg[39]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [39:36]),
        .S({\main_195_zSig0ii_reg[39]_i_6_n_0 ,\main_195_zSig0ii_reg[39]_i_7_n_0 ,\main_195_zSig0ii_reg[39]_i_8_n_0 ,\main_195_zSig0ii_reg[39]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\main_195_zSig0ii_reg_reg[3]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[3]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[3]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[3]_i_1_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\main_195_zSig0ii_reg[3]_i_2_n_0 ,\main_195_zSig0ii_reg[3]_i_3_n_0 ,\main_195_zSig0ii_reg[3]_i_4_n_0 ,\main_195_zSig0ii_reg[3]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [3:0]),
        .S({\main_195_zSig0ii_reg[3]_i_6_n_0 ,\main_195_zSig0ii_reg[3]_i_7_n_0 ,\main_195_zSig0ii_reg[3]_i_8_n_0 ,\main_195_zSig0ii_reg[3]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[43]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[39]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[43]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[43]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[43]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[43]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\main_195_zSig0ii_reg[43]_i_2_n_0 ,\main_195_zSig0ii_reg[43]_i_3_n_0 }),
        .O(\main_inst/main_195_zSig0ii [43:40]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\main_195_zSig0ii_reg[43]_i_4_n_0 ,\main_195_zSig0ii_reg[43]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[47]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[43]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[47]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[47]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[47]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[47]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O(\main_inst/main_195_zSig0ii [47:44]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[51]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[47]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[51]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[51]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[51]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[51]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O(\main_inst/main_195_zSig0ii [51:48]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[55]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[51]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[55]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[55]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[55]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[55]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O(\main_inst/main_195_zSig0ii [55:52]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[59]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[55]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[59]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[59]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[59]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[59]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O(\main_inst/main_195_zSig0ii [59:56]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[63]_i_2 
       (.CI(\main_195_zSig0ii_reg_reg[59]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O(\main_inst/main_195_zSig0ii [63:60]),
        .S({\<const1>__0__0 ,\main_195_zSig0ii_reg[63]_i_4_n_0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_195_zSig0ii_reg_reg[7]_i_1 
       (.CI(\main_195_zSig0ii_reg_reg[3]_i_1_n_0 ),
        .CO({\main_195_zSig0ii_reg_reg[7]_i_1_n_0 ,\main_195_zSig0ii_reg_reg[7]_i_1_n_1 ,\main_195_zSig0ii_reg_reg[7]_i_1_n_2 ,\main_195_zSig0ii_reg_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_195_zSig0ii_reg[7]_i_2_n_0 ,\main_195_zSig0ii_reg[7]_i_3_n_0 ,\main_195_zSig0ii_reg[7]_i_4_n_0 ,\main_195_zSig0ii_reg[7]_i_5_n_0 }),
        .O(\main_inst/main_195_zSig0ii [7:4]),
        .S({\main_195_zSig0ii_reg[7]_i_6_n_0 ,\main_195_zSig0ii_reg[7]_i_7_n_0 ,\main_195_zSig0ii_reg[7]_i_8_n_0 ,\main_195_zSig0ii_reg[7]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1000)) 
    \main_1_2_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .O(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000988810001000)) 
    \main_1_2_reg[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_float64_addexit_exitcond1_reg ),
        .I5(\main_1_2_reg[31]_i_4_n_0 ),
        .O(\main_inst/main_1_2_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \main_1_2_reg[31]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_1_2_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \main_1_2_reg[31]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_1_2_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \main_1_4_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(main_1_4_reg),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_inst/main_1_3_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_1_4_reg[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .O(main_1_4_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[0]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/CI ),
        .O(main_1_main_result02_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[0]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [3]),
        .O(\main_1_main_result02_reg[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[0]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [2]),
        .O(\main_1_main_result02_reg[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[0]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [1]),
        .O(\main_1_main_result02_reg[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000EFFFEFFF0000)) 
    \main_1_main_result02_reg[0]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/CI ),
        .I5(\main_inst/main_1_main_result02_reg_reg [0]),
        .O(\main_1_main_result02_reg[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[12]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [15]),
        .O(\main_1_main_result02_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[12]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [14]),
        .O(\main_1_main_result02_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[12]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [13]),
        .O(\main_1_main_result02_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[12]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [12]),
        .O(\main_1_main_result02_reg[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[16]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [19]),
        .O(\main_1_main_result02_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[16]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [18]),
        .O(\main_1_main_result02_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[16]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [17]),
        .O(\main_1_main_result02_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[16]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [16]),
        .O(\main_1_main_result02_reg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[20]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [23]),
        .O(\main_1_main_result02_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[20]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [22]),
        .O(\main_1_main_result02_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[20]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [21]),
        .O(\main_1_main_result02_reg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[20]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [20]),
        .O(\main_1_main_result02_reg[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[24]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [27]),
        .O(\main_1_main_result02_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[24]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [26]),
        .O(\main_1_main_result02_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[24]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [25]),
        .O(\main_1_main_result02_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[24]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [24]),
        .O(\main_1_main_result02_reg[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[28]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [31]),
        .O(\main_1_main_result02_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[28]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [30]),
        .O(\main_1_main_result02_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[28]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [29]),
        .O(\main_1_main_result02_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[28]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [28]),
        .O(\main_1_main_result02_reg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[4]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [7]),
        .O(\main_1_main_result02_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[4]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [6]),
        .O(\main_1_main_result02_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[4]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [5]),
        .O(\main_1_main_result02_reg[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[4]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [4]),
        .O(\main_1_main_result02_reg[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[8]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [11]),
        .O(\main_1_main_result02_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[8]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [10]),
        .O(\main_1_main_result02_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[8]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [9]),
        .O(\main_1_main_result02_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEFFF0000)) 
    \main_1_main_result02_reg[8]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_3_n_0 ),
        .I3(start),
        .I4(\main_inst/main_1_main_result02_reg_reg [8]),
        .O(\main_1_main_result02_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[0]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(main_1_main_result02_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,main_1_main_result02_reg}),
        .O({\main_1_main_result02_reg_reg[0]_i_1_n_4 ,\main_1_main_result02_reg_reg[0]_i_1_n_5 ,\main_1_main_result02_reg_reg[0]_i_1_n_6 ,\main_1_main_result02_reg_reg[0]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[0]_i_3_n_0 ,\main_1_main_result02_reg[0]_i_4_n_0 ,\main_1_main_result02_reg[0]_i_5_n_0 ,\main_1_main_result02_reg[0]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[12]_i_1 
       (.CI(\main_1_main_result02_reg_reg[8]_i_1_n_0 ),
        .CO({\main_1_main_result02_reg_reg[12]_i_1_n_0 ,\main_1_main_result02_reg_reg[12]_i_1_n_1 ,\main_1_main_result02_reg_reg[12]_i_1_n_2 ,\main_1_main_result02_reg_reg[12]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[12]_i_1_n_4 ,\main_1_main_result02_reg_reg[12]_i_1_n_5 ,\main_1_main_result02_reg_reg[12]_i_1_n_6 ,\main_1_main_result02_reg_reg[12]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[12]_i_2_n_0 ,\main_1_main_result02_reg[12]_i_3_n_0 ,\main_1_main_result02_reg[12]_i_4_n_0 ,\main_1_main_result02_reg[12]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[16]_i_1 
       (.CI(\main_1_main_result02_reg_reg[12]_i_1_n_0 ),
        .CO({\main_1_main_result02_reg_reg[16]_i_1_n_0 ,\main_1_main_result02_reg_reg[16]_i_1_n_1 ,\main_1_main_result02_reg_reg[16]_i_1_n_2 ,\main_1_main_result02_reg_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[16]_i_1_n_4 ,\main_1_main_result02_reg_reg[16]_i_1_n_5 ,\main_1_main_result02_reg_reg[16]_i_1_n_6 ,\main_1_main_result02_reg_reg[16]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[16]_i_2_n_0 ,\main_1_main_result02_reg[16]_i_3_n_0 ,\main_1_main_result02_reg[16]_i_4_n_0 ,\main_1_main_result02_reg[16]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[20]_i_1 
       (.CI(\main_1_main_result02_reg_reg[16]_i_1_n_0 ),
        .CO({\main_1_main_result02_reg_reg[20]_i_1_n_0 ,\main_1_main_result02_reg_reg[20]_i_1_n_1 ,\main_1_main_result02_reg_reg[20]_i_1_n_2 ,\main_1_main_result02_reg_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[20]_i_1_n_4 ,\main_1_main_result02_reg_reg[20]_i_1_n_5 ,\main_1_main_result02_reg_reg[20]_i_1_n_6 ,\main_1_main_result02_reg_reg[20]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[20]_i_2_n_0 ,\main_1_main_result02_reg[20]_i_3_n_0 ,\main_1_main_result02_reg[20]_i_4_n_0 ,\main_1_main_result02_reg[20]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[24]_i_1 
       (.CI(\main_1_main_result02_reg_reg[20]_i_1_n_0 ),
        .CO({\main_1_main_result02_reg_reg[24]_i_1_n_0 ,\main_1_main_result02_reg_reg[24]_i_1_n_1 ,\main_1_main_result02_reg_reg[24]_i_1_n_2 ,\main_1_main_result02_reg_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[24]_i_1_n_4 ,\main_1_main_result02_reg_reg[24]_i_1_n_5 ,\main_1_main_result02_reg_reg[24]_i_1_n_6 ,\main_1_main_result02_reg_reg[24]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[24]_i_2_n_0 ,\main_1_main_result02_reg[24]_i_3_n_0 ,\main_1_main_result02_reg[24]_i_4_n_0 ,\main_1_main_result02_reg[24]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[28]_i_1 
       (.CI(\main_1_main_result02_reg_reg[24]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[28]_i_1_n_4 ,\main_1_main_result02_reg_reg[28]_i_1_n_5 ,\main_1_main_result02_reg_reg[28]_i_1_n_6 ,\main_1_main_result02_reg_reg[28]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[28]_i_2_n_0 ,\main_1_main_result02_reg[28]_i_3_n_0 ,\main_1_main_result02_reg[28]_i_4_n_0 ,\main_1_main_result02_reg[28]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[4]_i_1 
       (.CI(main_1_main_result02_reg_reg[3]),
        .CO({\main_1_main_result02_reg_reg[4]_i_1_n_0 ,\main_1_main_result02_reg_reg[4]_i_1_n_1 ,\main_1_main_result02_reg_reg[4]_i_1_n_2 ,\main_1_main_result02_reg_reg[4]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[4]_i_1_n_4 ,\main_1_main_result02_reg_reg[4]_i_1_n_5 ,\main_1_main_result02_reg_reg[4]_i_1_n_6 ,\main_1_main_result02_reg_reg[4]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[4]_i_2_n_0 ,\main_1_main_result02_reg[4]_i_3_n_0 ,\main_1_main_result02_reg[4]_i_4_n_0 ,\main_1_main_result02_reg[4]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_main_result02_reg_reg[8]_i_1 
       (.CI(\main_1_main_result02_reg_reg[4]_i_1_n_0 ),
        .CO({\main_1_main_result02_reg_reg[8]_i_1_n_0 ,\main_1_main_result02_reg_reg[8]_i_1_n_1 ,\main_1_main_result02_reg_reg[8]_i_1_n_2 ,\main_1_main_result02_reg_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_main_result02_reg_reg[8]_i_1_n_4 ,\main_1_main_result02_reg_reg[8]_i_1_n_5 ,\main_1_main_result02_reg_reg[8]_i_1_n_6 ,\main_1_main_result02_reg_reg[8]_i_1_n_7 }),
        .S({\main_1_main_result02_reg[8]_i_2_n_0 ,\main_1_main_result02_reg[8]_i_3_n_0 ,\main_1_main_result02_reg[8]_i_4_n_0 ,\main_1_main_result02_reg[8]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \main_1_scevgep_reg[25]_i_2 
       (.I0(\main_inst/main_1_scevgep_reg1 [25]),
        .O(main_1_scevgep_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \main_1_scevgep_reg[25]_i_4 
       (.I0(\main_inst/main_1_scevgep_reg1 [23]),
        .O(\main_1_scevgep_reg[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \main_1_scevgep_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_1_scevgep_reg[31]_i_3_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_inst/main_1_scevgep_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_1_scevgep_reg[31]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_1_scevgep_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_scevgep_reg_reg[25]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(main_1_scevgep_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_1_scevgep_reg1 [25],\<const0>__0__0 ,\main_inst/main_1_scevgep_reg1 [23],\<const0>__0__0 }),
        .O({\main_inst/main_1_scevgep [25:23],\main_1_scevgep_reg_reg[25]_i_1_n_7 }),
        .S({main_1_scevgep_reg,\main_inst/main_1_scevgep_reg1 [24],\main_1_scevgep_reg[25]_i_4_n_0 ,\main_inst/main_1_scevgep_reg1 [22]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_scevgep_reg_reg[29]_i_1 
       (.CI(main_1_scevgep_reg_reg[3]),
        .CO({\main_1_scevgep_reg_reg[29]_i_1_n_0 ,\main_1_scevgep_reg_reg[29]_i_1_n_1 ,\main_1_scevgep_reg_reg[29]_i_1_n_2 ,\main_1_scevgep_reg_reg[29]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_1_scevgep [29:26]),
        .S(\main_inst/main_1_scevgep_reg1 [29:26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_1_scevgep_reg_reg[31]_i_2 
       (.CI(\main_1_scevgep_reg_reg[29]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_1_scevgep_reg_reg[31]_i_2_n_4 ,\main_1_scevgep_reg_reg[31]_i_2_n_5 ,\main_inst/main_1_scevgep [31:30]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_1_scevgep_reg1 [31:30]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000004)) 
    \main_27_expDiff0i2i_reg[31]_i_1 
       (.I0(main_27_expDiff0i2i_reg),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_inst/main_27_30_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFD)) 
    \main_27_expDiff0i2i_reg[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .O(main_27_expDiff0i2i_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000040)) 
    \main_59_expDiff1i3i_reg[31]_i_1 
       (.I0(main_27_expDiff0i2i_reg),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_inst/main_59_62_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[0]_i_1 
       (.I0(\main_float64_addexit_0i_reg[0]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[0]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[0]_i_4_n_0 ),
        .O(main_float64_addexit_0i_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[0]_i_2 
       (.I0(\main_float64_addexit_0i_reg[0]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [9]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[0]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_ ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [9]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[0]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[0]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [9]),
        .O(\main_float64_addexit_0i_reg[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[0]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_ ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [9]),
        .O(\main_float64_addexit_0i_reg[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAA3CAA00)) 
    \main_float64_addexit_0i_reg[0]_i_6 
       (.I0(\main_inst/main_15_17 [9]),
        .I1(\main_inst/main_15_19_reg [9]),
        .I2(\main_inst/main_91_92 [9]),
        .I3(\main_inst/main_float64_addexit_0i121_out ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[10]_i_1 
       (.I0(\main_float64_addexit_0i_reg[10]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[10]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[10]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[10]_i_2 
       (.I0(\main_float64_addexit_0i_reg[10]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [19]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[10]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[10] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [19]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[10]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[10]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [19]),
        .O(\main_float64_addexit_0i_reg[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[10]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[10] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [19]),
        .O(\main_float64_addexit_0i_reg[10]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[10]_i_6 
       (.I0(\main_inst/main_15_17 [19]),
        .I1(\main_inst/data5 [10]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[10]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[11]_i_1 
       (.I0(\main_float64_addexit_0i_reg[11]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[11]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[11]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[11]_i_10 
       (.I0(\main_inst/main_15_19_reg [18]),
        .I1(\main_inst/main_91_92 [18]),
        .O(\main_float64_addexit_0i_reg[11]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[11]_i_11 
       (.I0(\main_inst/main_15_19_reg [17]),
        .I1(\main_inst/main_91_92 [17]),
        .O(\main_float64_addexit_0i_reg[11]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[11]_i_2 
       (.I0(\main_float64_addexit_0i_reg[11]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [20]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[11]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[11] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [20]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[11]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[11]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [20]),
        .O(\main_float64_addexit_0i_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[11]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[11] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [20]),
        .O(\main_float64_addexit_0i_reg[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[11]_i_6 
       (.I0(\main_inst/main_15_17 [20]),
        .I1(\main_inst/data5 [11]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[11]_i_8 
       (.I0(\main_inst/main_15_19_reg [20]),
        .I1(\main_inst/main_91_92 [20]),
        .O(\main_float64_addexit_0i_reg[11]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[11]_i_9 
       (.I0(\main_inst/main_15_19_reg [19]),
        .I1(\main_inst/main_91_92 [19]),
        .O(\main_float64_addexit_0i_reg[11]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[12]_i_1 
       (.I0(\main_float64_addexit_0i_reg[12]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[12]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[12]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[12]_i_2 
       (.I0(\main_float64_addexit_0i_reg[12]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [21]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[12]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[12] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [21]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[12]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[12]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [21]),
        .O(\main_float64_addexit_0i_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[12]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[12] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [21]),
        .O(\main_float64_addexit_0i_reg[12]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[12]_i_6 
       (.I0(\main_inst/main_15_17 [21]),
        .I1(\main_inst/data5 [12]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[12]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[13]_i_1 
       (.I0(\main_float64_addexit_0i_reg[13]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[13]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[13]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[13]_i_2 
       (.I0(\main_float64_addexit_0i_reg[13]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [22]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[13]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[13] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [22]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[13]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[13]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [22]),
        .O(\main_float64_addexit_0i_reg[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[13]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [22]),
        .O(\main_float64_addexit_0i_reg[13]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[13]_i_6 
       (.I0(\main_inst/main_15_17 [22]),
        .I1(\main_inst/data5 [13]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[13]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[14]_i_1 
       (.I0(\main_float64_addexit_0i_reg[14]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[14]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[14]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[14]_i_2 
       (.I0(\main_float64_addexit_0i_reg[14]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [23]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[14]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[14] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [23]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[14]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[14]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [23]),
        .O(\main_float64_addexit_0i_reg[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[14]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [23]),
        .O(\main_float64_addexit_0i_reg[14]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[14]_i_6 
       (.I0(\main_inst/main_15_17 [23]),
        .I1(\main_inst/data5 [14]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[14]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[15]_i_1 
       (.I0(\main_float64_addexit_0i_reg[15]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[15]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[15]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[15]_i_10 
       (.I0(\main_inst/main_15_19_reg [22]),
        .I1(\main_inst/main_91_92 [22]),
        .O(\main_float64_addexit_0i_reg[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[15]_i_11 
       (.I0(\main_inst/main_15_19_reg [21]),
        .I1(\main_inst/main_91_92 [21]),
        .O(\main_float64_addexit_0i_reg[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[15]_i_2 
       (.I0(\main_float64_addexit_0i_reg[15]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [24]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[15]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[15] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [24]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[15]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[15]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [24]),
        .O(\main_float64_addexit_0i_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[15]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[15] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [24]),
        .O(\main_float64_addexit_0i_reg[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[15]_i_6 
       (.I0(\main_inst/main_15_17 [24]),
        .I1(\main_inst/data5 [15]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[15]_i_8 
       (.I0(\main_inst/main_15_19_reg [24]),
        .I1(\main_inst/main_91_92 [24]),
        .O(\main_float64_addexit_0i_reg[15]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[15]_i_9 
       (.I0(\main_inst/main_15_19_reg [23]),
        .I1(\main_inst/main_91_92 [23]),
        .O(\main_float64_addexit_0i_reg[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[16]_i_1 
       (.I0(\main_float64_addexit_0i_reg[16]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[16]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[16]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[16]_i_2 
       (.I0(\main_float64_addexit_0i_reg[16]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [25]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[16]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[16] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [25]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[16]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[16]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [25]),
        .O(\main_float64_addexit_0i_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[16]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [25]),
        .O(\main_float64_addexit_0i_reg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[16]_i_6 
       (.I0(\main_inst/main_15_17 [25]),
        .I1(\main_inst/data5 [16]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[17]_i_1 
       (.I0(\main_float64_addexit_0i_reg[17]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[17]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[17]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[17]_i_2 
       (.I0(\main_float64_addexit_0i_reg[17]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [26]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[17]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[17] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [26]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[17]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[17]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [26]),
        .O(\main_float64_addexit_0i_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[17]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[17] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [26]),
        .O(\main_float64_addexit_0i_reg[17]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[17]_i_6 
       (.I0(\main_inst/main_15_17 [26]),
        .I1(\main_inst/data5 [17]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[17]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[18]_i_1 
       (.I0(\main_float64_addexit_0i_reg[18]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[18]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[18]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[18]_i_2 
       (.I0(\main_float64_addexit_0i_reg[18]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [27]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[18]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[18] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [27]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[18]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[18]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [27]),
        .O(\main_float64_addexit_0i_reg[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[18]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[18] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [27]),
        .O(\main_float64_addexit_0i_reg[18]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[18]_i_6 
       (.I0(\main_inst/main_15_17 [27]),
        .I1(\main_inst/data5 [18]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[18]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[19]_i_1 
       (.I0(\main_float64_addexit_0i_reg[19]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[19]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[19]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[19]_i_10 
       (.I0(\main_inst/main_15_19_reg [26]),
        .I1(\main_inst/main_91_92 [26]),
        .O(\main_float64_addexit_0i_reg[19]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[19]_i_11 
       (.I0(\main_inst/main_15_19_reg [25]),
        .I1(\main_inst/main_91_92 [25]),
        .O(\main_float64_addexit_0i_reg[19]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[19]_i_2 
       (.I0(\main_float64_addexit_0i_reg[19]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [28]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[19]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[19] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [28]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[19]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[19]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [28]),
        .O(\main_float64_addexit_0i_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[19]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [28]),
        .O(\main_float64_addexit_0i_reg[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[19]_i_6 
       (.I0(\main_inst/main_15_17 [28]),
        .I1(\main_inst/data5 [19]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[19]_i_8 
       (.I0(\main_inst/main_15_19_reg [28]),
        .I1(\main_inst/main_91_92 [28]),
        .O(\main_float64_addexit_0i_reg[19]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[19]_i_9 
       (.I0(\main_inst/main_15_19_reg [27]),
        .I1(\main_inst/main_91_92 [27]),
        .O(\main_float64_addexit_0i_reg[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[1]_i_1 
       (.I0(\main_float64_addexit_0i_reg[1]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[1]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[1]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[1]_i_2 
       (.I0(\main_float64_addexit_0i_reg[1]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [10]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[1]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[1] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [10]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[1]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[1]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [10]),
        .O(\main_float64_addexit_0i_reg[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[1]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[1] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [10]),
        .O(\main_float64_addexit_0i_reg[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[1]_i_6 
       (.I0(\main_inst/main_15_17 [10]),
        .I1(\main_inst/data5 [1]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[1]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[20]_i_1 
       (.I0(\main_float64_addexit_0i_reg[20]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[20]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[20]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[20]_i_2 
       (.I0(\main_float64_addexit_0i_reg[20]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [29]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[20]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[20] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [29]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[20]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[20]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [29]),
        .O(\main_float64_addexit_0i_reg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[20]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [29]),
        .O(\main_float64_addexit_0i_reg[20]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[20]_i_6 
       (.I0(\main_inst/main_15_17 [29]),
        .I1(\main_inst/data5 [20]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[20]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[21]_i_1 
       (.I0(\main_float64_addexit_0i_reg[21]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[21]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[21]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[21]_i_2 
       (.I0(\main_float64_addexit_0i_reg[21]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [30]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[21]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[21] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [30]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[21]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[21]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [30]),
        .O(\main_float64_addexit_0i_reg[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[21]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[21] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [30]),
        .O(\main_float64_addexit_0i_reg[21]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[21]_i_6 
       (.I0(\main_inst/main_15_17 [30]),
        .I1(\main_inst/data5 [21]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[21]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[22]_i_1 
       (.I0(\main_float64_addexit_0i_reg[22]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[22]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[22]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[22]_i_2 
       (.I0(\main_float64_addexit_0i_reg[22]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [31]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[22]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[22] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [31]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[22]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[22]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [31]),
        .O(\main_float64_addexit_0i_reg[22]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[22]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [31]),
        .O(\main_float64_addexit_0i_reg[22]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[22]_i_6 
       (.I0(\main_inst/main_15_17 [31]),
        .I1(\main_inst/data5 [22]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[22]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[23]_i_1 
       (.I0(\main_float64_addexit_0i_reg[23]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[23]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[23]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[23]_i_10 
       (.I0(\main_inst/main_15_19_reg [30]),
        .I1(\main_inst/main_91_92 [30]),
        .O(\main_float64_addexit_0i_reg[23]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[23]_i_11 
       (.I0(\main_inst/main_15_19_reg [29]),
        .I1(\main_inst/main_91_92 [29]),
        .O(\main_float64_addexit_0i_reg[23]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[23]_i_2 
       (.I0(\main_float64_addexit_0i_reg[23]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [32]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[23]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[23] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [32]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[23]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[23]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [32]),
        .O(\main_float64_addexit_0i_reg[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[23]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[23] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [32]),
        .O(\main_float64_addexit_0i_reg[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[23]_i_6 
       (.I0(\main_inst/main_15_17 [32]),
        .I1(\main_inst/data5 [23]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[23]_i_8 
       (.I0(\main_inst/main_15_19_reg [32]),
        .I1(\main_inst/main_91_92 [32]),
        .O(\main_float64_addexit_0i_reg[23]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[23]_i_9 
       (.I0(\main_inst/main_15_19_reg [31]),
        .I1(\main_inst/main_91_92 [31]),
        .O(\main_float64_addexit_0i_reg[23]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[24]_i_1 
       (.I0(\main_float64_addexit_0i_reg[24]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[24]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[24]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[24]_i_2 
       (.I0(\main_float64_addexit_0i_reg[24]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [33]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[24]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[24] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [33]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[24]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[24]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [33]),
        .O(\main_float64_addexit_0i_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[24]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[24] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [33]),
        .O(\main_float64_addexit_0i_reg[24]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[24]_i_6 
       (.I0(\main_inst/main_15_17 [33]),
        .I1(\main_inst/data5 [24]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[24]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[25]_i_1 
       (.I0(\main_float64_addexit_0i_reg[25]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[25]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[25]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[25]_i_2 
       (.I0(\main_float64_addexit_0i_reg[25]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [34]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[25]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[25] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [34]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[25]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[25]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [34]),
        .O(\main_float64_addexit_0i_reg[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[25]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [34]),
        .O(\main_float64_addexit_0i_reg[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[25]_i_6 
       (.I0(\main_inst/main_15_17 [34]),
        .I1(\main_inst/data5 [25]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[25]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[26]_i_1 
       (.I0(\main_float64_addexit_0i_reg[26]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[26]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[26]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[26]_i_2 
       (.I0(\main_float64_addexit_0i_reg[26]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [35]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[26]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[26] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [35]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[26]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[26]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [35]),
        .O(\main_float64_addexit_0i_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[26]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [35]),
        .O(\main_float64_addexit_0i_reg[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[26]_i_6 
       (.I0(\main_inst/main_15_17 [35]),
        .I1(\main_inst/data5 [26]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[26]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[27]_i_1 
       (.I0(\main_float64_addexit_0i_reg[27]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[27]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[27]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[27]_i_2 
       (.I0(\main_float64_addexit_0i_reg[27]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [36]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[27]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[27] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [36]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[27]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[27]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [36]),
        .O(\main_float64_addexit_0i_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[27]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[27] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [36]),
        .O(\main_float64_addexit_0i_reg[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[27]_i_6 
       (.I0(\main_inst/main_15_17 [36]),
        .I1(\main_inst/data5 [27]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[28]_i_1 
       (.I0(\main_float64_addexit_0i_reg[28]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[28]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[28]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[28]_i_2 
       (.I0(\main_float64_addexit_0i_reg[28]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [37]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[28]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[28] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [37]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[28]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[28]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [37]),
        .O(\main_float64_addexit_0i_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[28]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [37]),
        .O(\main_float64_addexit_0i_reg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[28]_i_6 
       (.I0(\main_inst/main_15_17 [37]),
        .I1(\main_inst/data5 [28]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[28]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[29]_i_1 
       (.I0(\main_float64_addexit_0i_reg[29]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[29]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[29]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[29]_i_2 
       (.I0(\main_float64_addexit_0i_reg[29]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [38]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[29]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[29] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [38]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[29]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[29]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [38]),
        .O(\main_float64_addexit_0i_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[29]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[29] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [38]),
        .O(\main_float64_addexit_0i_reg[29]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[29]_i_6 
       (.I0(\main_inst/main_15_17 [38]),
        .I1(\main_inst/data5 [29]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[29]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[2]_i_1 
       (.I0(\main_float64_addexit_0i_reg[2]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[2]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[2]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[2]_i_2 
       (.I0(\main_float64_addexit_0i_reg[2]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [11]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[2]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[2] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [11]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[2]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[2]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [11]),
        .O(\main_float64_addexit_0i_reg[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[2]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[2] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [11]),
        .O(\main_float64_addexit_0i_reg[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[2]_i_6 
       (.I0(\main_inst/main_15_17 [11]),
        .I1(\main_inst/data5 [2]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[30]_i_1 
       (.I0(\main_float64_addexit_0i_reg[30]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[30]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[30]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[30]_i_2 
       (.I0(\main_float64_addexit_0i_reg[30]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [39]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[30]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[30] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [39]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[30]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[30]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [39]),
        .O(\main_float64_addexit_0i_reg[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[30]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[30] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [39]),
        .O(\main_float64_addexit_0i_reg[30]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[30]_i_6 
       (.I0(\main_inst/main_15_17 [39]),
        .I1(\main_inst/data5 [30]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[30]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[31]_i_1 
       (.I0(\main_float64_addexit_0i_reg[31]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[31]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[31]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[31]_i_2 
       (.I0(\main_float64_addexit_0i_reg[31]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [40]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[31]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[31] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [40]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[31]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[31]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [40]),
        .O(\main_float64_addexit_0i_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[31]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [40]),
        .O(\main_float64_addexit_0i_reg[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[31]_i_6 
       (.I0(\main_inst/main_15_17 [40]),
        .I1(\main_inst/data5 [31]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'hF4)) 
    \main_float64_addexit_0i_reg[32]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[32]_i_2_n_0 ),
        .I2(\main_float64_addexit_0i_reg[32]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_10 
       (.I0(\main_inst/main_15_19_reg [37]),
        .I1(\main_inst/main_91_92 [37]),
        .O(\main_float64_addexit_0i_reg[32]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_11 
       (.I0(\main_inst/main_15_19_reg [36]),
        .I1(\main_inst/main_91_92 [36]),
        .O(\main_float64_addexit_0i_reg[32]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_12 
       (.I0(\main_inst/main_15_19_reg [35]),
        .I1(\main_inst/main_91_92 [35]),
        .O(\main_float64_addexit_0i_reg[32]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_13 
       (.I0(\main_inst/main_15_19_reg [34]),
        .I1(\main_inst/main_91_92 [34]),
        .O(\main_float64_addexit_0i_reg[32]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_14 
       (.I0(\main_inst/main_15_19_reg [33]),
        .I1(\main_inst/main_91_92 [33]),
        .O(\main_float64_addexit_0i_reg[32]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[32]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[32] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[32]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \main_float64_addexit_0i_reg[32]_i_3 
       (.I0(\main_inst/data5 [32]),
        .I1(\main_inst/main_float64_addexit_0i129_out ),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .O(\main_float64_addexit_0i_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[32]_i_4 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[32] ),
        .O(\main_float64_addexit_0i_reg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_7 
       (.I0(\main_inst/main_15_19_reg [40]),
        .I1(\main_inst/main_91_92 [40]),
        .O(\main_float64_addexit_0i_reg[32]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_8 
       (.I0(\main_inst/main_15_19_reg [39]),
        .I1(\main_inst/main_91_92 [39]),
        .O(\main_float64_addexit_0i_reg[32]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[32]_i_9 
       (.I0(\main_inst/main_15_19_reg [38]),
        .I1(\main_inst/main_91_92 [38]),
        .O(\main_float64_addexit_0i_reg[32]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[33]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[33]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[33]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[33] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[33]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[33]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[33] ),
        .O(\main_float64_addexit_0i_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[34]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[34]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[34]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[34]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[34] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[34]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[34]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[34] ),
        .O(\main_float64_addexit_0i_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[35]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[35]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[35]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[35]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[35] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[35]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[35]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[35] ),
        .O(\main_float64_addexit_0i_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[36]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[36]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[36]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[36]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[36] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[36]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[36]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[36] ),
        .O(\main_float64_addexit_0i_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[37]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[37]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[37]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[37]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[37] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[37]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[37]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[37] ),
        .O(\main_float64_addexit_0i_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[38]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[38]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[38]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[38]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[38] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[38]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[38]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[38] ),
        .O(\main_float64_addexit_0i_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[39]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[39]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[39]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[39]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[39] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[39]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[39]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[39] ),
        .O(\main_float64_addexit_0i_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[3]_i_1 
       (.I0(\main_float64_addexit_0i_reg[3]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[3]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[3]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[3]_i_10 
       (.I0(\main_inst/main_15_19_reg [10]),
        .I1(\main_inst/main_91_92 [10]),
        .O(\main_float64_addexit_0i_reg[3]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[3]_i_11 
       (.I0(\main_inst/main_15_19_reg [9]),
        .I1(\main_inst/main_91_92 [9]),
        .O(\main_inst/data5 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[3]_i_2 
       (.I0(\main_float64_addexit_0i_reg[3]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [12]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[3]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[3] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [12]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[3]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[3]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [12]),
        .O(\main_float64_addexit_0i_reg[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[3]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[3] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [12]),
        .O(\main_float64_addexit_0i_reg[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[3]_i_6 
       (.I0(\main_inst/main_15_17 [12]),
        .I1(\main_inst/data5 [3]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[3]_i_8 
       (.I0(\main_inst/main_15_19_reg [12]),
        .I1(\main_inst/main_91_92 [12]),
        .O(\main_float64_addexit_0i_reg[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[3]_i_9 
       (.I0(\main_inst/main_15_19_reg [11]),
        .I1(\main_inst/main_91_92 [11]),
        .O(\main_float64_addexit_0i_reg[3]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[40]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[40]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[40]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[40]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[40] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[40]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[40]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[40] ),
        .O(\main_float64_addexit_0i_reg[40]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[41]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[41]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[41]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[41] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[41]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[41]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[41]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[41] ),
        .O(\main_float64_addexit_0i_reg[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[42]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[42]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[42]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[42]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[42] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[42]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[42]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[42]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[42] ),
        .O(\main_float64_addexit_0i_reg[42]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[43]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[43]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[43]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[43]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[43] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[43]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[43]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[43]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[43] ),
        .O(\main_float64_addexit_0i_reg[43]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[44]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[44]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[44]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[44]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[44] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[44]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[44]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[44]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[44] ),
        .O(\main_float64_addexit_0i_reg[44]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[45]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[45]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[45]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[45]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[45] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[45]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[45]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[45]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[45] ),
        .O(\main_float64_addexit_0i_reg[45]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[46]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[46]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[46]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[46]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[46] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[46]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[46]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[46]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[46] ),
        .O(\main_float64_addexit_0i_reg[46]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[47]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[47]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[47]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[47]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[47] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[47]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[47]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[47]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[47] ),
        .O(\main_float64_addexit_0i_reg[47]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[48]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[48]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[48]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[48]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[48] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[48]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[48]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[48]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[48] ),
        .O(\main_float64_addexit_0i_reg[48]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[49]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[49]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[49]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[49]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[49] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[49]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[49]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[49] ),
        .O(\main_float64_addexit_0i_reg[49]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[4]_i_1 
       (.I0(\main_float64_addexit_0i_reg[4]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[4]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[4]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[4]_i_2 
       (.I0(\main_float64_addexit_0i_reg[4]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [13]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[4]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[4] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [13]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[4]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[4]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [13]),
        .O(\main_float64_addexit_0i_reg[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[4]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[4] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [13]),
        .O(\main_float64_addexit_0i_reg[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[4]_i_6 
       (.I0(\main_inst/main_15_17 [13]),
        .I1(\main_inst/data5 [4]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT2 #(
    .INIT(4'h4)) 
    \main_float64_addexit_0i_reg[50]_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I1(\main_float64_addexit_0i_reg[50]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[50]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000400000004)) 
    \main_float64_addexit_0i_reg[50]_i_2 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[50] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[50]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[50]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \main_float64_addexit_0i_reg[50]_i_3 
       (.I0(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_inst/main_101_102_reg_reg_n_0_[50] ),
        .O(\main_float64_addexit_0i_reg[50]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \main_float64_addexit_0i_reg[51]_i_1 
       (.I0(\main_float64_addexit_0i_reg[51]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I2(\main_float64_addexit_0i_reg[51]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[51]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF5D0800005D08)) 
    \main_float64_addexit_0i_reg[51]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_float64_addexit_0i_reg[51]_i_4_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I5(\main_float64_addexit_0i_reg[51]_i_5_n_0 ),
        .O(\main_float64_addexit_0i_reg[51]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0F0F0F0004040404)) 
    \main_float64_addexit_0i_reg[51]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i121_out ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .I2(\main_inst/main_float64_addexit_0i129_out ),
        .I3(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I4(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .O(\main_float64_addexit_0i_reg[51]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h32)) 
    \main_float64_addexit_0i_reg[51]_i_4 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[51] ),
        .I1(\main_inst/main_float64_addexit_0i13_out ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .O(\main_float64_addexit_0i_reg[51]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFECE)) 
    \main_float64_addexit_0i_reg[51]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I3(\main_inst/main_101_102_reg_reg_n_0_[51] ),
        .O(\main_float64_addexit_0i_reg[51]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE2)) 
    \main_float64_addexit_0i_reg[52]_i_1 
       (.I0(\main_float64_addexit_0i_reg[52]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I2(\main_float64_addexit_0i_reg[52]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[52]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[52]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[52]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[52] ),
        .O(\main_float64_addexit_0i_reg[52]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[52]_i_4 
       (.I0(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_inst/main_float64_addexit_0i129_out ),
        .O(\main_float64_addexit_0i_reg[52]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[52]_i_5 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[52] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[52]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[53]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[53]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[53]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[53]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[53]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[53] ),
        .O(\main_float64_addexit_0i_reg[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[53]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[53] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[53]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[54]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[54]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[54]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[54]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[54]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[54] ),
        .O(\main_float64_addexit_0i_reg[54]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[54]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[54] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[54]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[55]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[55]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[55]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[55]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[55]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[55] ),
        .O(\main_float64_addexit_0i_reg[55]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[55]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[55] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[55]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[56]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[56]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[56]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[56]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[56]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[56] ),
        .O(\main_float64_addexit_0i_reg[56]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[56]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[56] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[56]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[57]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[57]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[57]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[57]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[57]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[57] ),
        .O(\main_float64_addexit_0i_reg[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[57]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[57] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[58]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[58]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[58]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[58]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[58]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[58] ),
        .O(\main_float64_addexit_0i_reg[58]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[58]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[58] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[58]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[59]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[59]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[59]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[59]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[59]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[59] ),
        .O(\main_float64_addexit_0i_reg[59]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[59]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[59] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[59]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[5]_i_1 
       (.I0(\main_float64_addexit_0i_reg[5]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[5]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[5]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[5]_i_2 
       (.I0(\main_float64_addexit_0i_reg[5]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [14]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[5]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[5] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [14]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[5]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[5]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [14]),
        .O(\main_float64_addexit_0i_reg[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[5]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[5] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [14]),
        .O(\main_float64_addexit_0i_reg[5]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[5]_i_6 
       (.I0(\main_inst/main_15_17 [14]),
        .I1(\main_inst/data5 [5]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[5]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[60]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[60]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[60]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[60]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[60]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[60] ),
        .O(\main_float64_addexit_0i_reg[60]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[60]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[60] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[60]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[61]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[61]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[61]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[61]_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[61]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[61] ),
        .O(\main_float64_addexit_0i_reg[61]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[61]_i_3 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[61] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[61]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \main_float64_addexit_0i_reg[62]_i_1 
       (.I0(\main_inst/main_float64_addexit_0i129_out ),
        .I1(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I5(\main_float64_addexit_0i_reg[62]_i_6_n_0 ),
        .O(\main_float64_addexit_0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000010000000)) 
    \main_float64_addexit_0i_reg[62]_i_10 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_158_160_reg[62]_i_4_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_float64_addexit_0i_reg[62]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_float64_addexit_0i_reg[62]_i_14 
       (.I0(\main_inst/main_91_92 [40]),
        .I1(\main_inst/main_91_92 [39]),
        .O(\main_float64_addexit_0i_reg[62]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_15 
       (.I0(\main_inst/main_91_92 [38]),
        .I1(\main_inst/main_91_92 [37]),
        .I2(\main_inst/main_91_92 [36]),
        .O(\main_float64_addexit_0i_reg[62]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_16 
       (.I0(\main_inst/main_91_92 [35]),
        .I1(\main_inst/main_91_92 [34]),
        .I2(\main_inst/main_91_92 [33]),
        .O(\main_float64_addexit_0i_reg[62]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_18 
       (.I0(\main_inst/main_91_92 [32]),
        .I1(\main_inst/main_91_92 [31]),
        .I2(\main_inst/main_91_92 [30]),
        .O(\main_float64_addexit_0i_reg[62]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_19 
       (.I0(\main_inst/main_91_92 [29]),
        .I1(\main_inst/main_91_92 [28]),
        .I2(\main_inst/main_91_92 [27]),
        .O(\main_float64_addexit_0i_reg[62]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \main_float64_addexit_0i_reg[62]_i_2 
       (.I0(\main_inst/main_23_24 ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_101_zExp1ii_reg[31]_i_3_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_inst/main_float64_addexit_0i129_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_20 
       (.I0(\main_inst/main_91_92 [26]),
        .I1(\main_inst/main_91_92 [25]),
        .I2(\main_inst/main_91_92 [24]),
        .O(\main_float64_addexit_0i_reg[62]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_21 
       (.I0(\main_inst/main_91_92 [23]),
        .I1(\main_inst/main_91_92 [22]),
        .I2(\main_inst/main_91_92 [21]),
        .O(\main_float64_addexit_0i_reg[62]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_22 
       (.I0(\main_inst/main_91_92 [20]),
        .I1(\main_inst/main_91_92 [19]),
        .I2(\main_inst/main_91_92 [18]),
        .O(\main_float64_addexit_0i_reg[62]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_23 
       (.I0(\main_inst/main_91_92 [17]),
        .I1(\main_inst/main_91_92 [16]),
        .I2(\main_inst/main_91_92 [15]),
        .O(\main_float64_addexit_0i_reg[62]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_24 
       (.I0(\main_inst/main_91_92 [14]),
        .I1(\main_inst/main_91_92 [13]),
        .I2(\main_inst/main_91_92 [12]),
        .O(\main_float64_addexit_0i_reg[62]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_0i_reg[62]_i_25 
       (.I0(\main_inst/main_91_92 [11]),
        .I1(\main_inst/main_91_92 [10]),
        .I2(\main_inst/main_91_92 [9]),
        .O(\main_float64_addexit_0i_reg[62]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    \main_float64_addexit_0i_reg[62]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(main_158_160_reg),
        .O(\main_float64_addexit_0i_reg[62]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \main_float64_addexit_0i_reg[62]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[62]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_float64_addexit_0i_reg[62]_i_5 
       (.I0(\main_float64_addexit_0i_reg[62]_i_8_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_float64_addexit_0i_reg[62]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFEFEAEFEAEFEAE)) 
    \main_float64_addexit_0i_reg[62]_i_6 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I5(\main_inst/main_101_102_reg_reg_n_0_[62] ),
        .O(\main_float64_addexit_0i_reg[62]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \main_float64_addexit_0i_reg[62]_i_8 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_float64_addexit_0i_reg[62]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[62]_i_9 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[62] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[62]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_1 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_3_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_4_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .O(\main_inst/main_float64_addexit_0i_reg0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_float64_addexit_0i_reg[63]_inv_i_10 
       (.I0(\main_inst/main_float64_addexit_0i13_out ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[63] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000004)) 
    \main_float64_addexit_0i_reg[63]_inv_i_11 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_23_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFFE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_12 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0800000000000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_13 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_158_160_reg[62]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_14 
       (.I0(\main_inst/main_165_166 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .O(\main_inst/main_float64_addexit_0i13_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00000400)) 
    \main_float64_addexit_0i_reg[63]_inv_i_15 
       (.I0(main_158_160_reg),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_inst/main_float64_addexit_0i129_out ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000008000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_16 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .I3(\main_inst/cur_state_reg_n_0_ ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/main_123_124 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000002000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_17 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_158_160_reg[62]_i_4_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0100400000000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_18 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_158_160_reg[62]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \main_float64_addexit_0i_reg[63]_inv_i_19 
       (.I0(\main_inst/main_81_83 ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_20_n_0 ),
        .O(\main_inst/main_float64_addexit_0i121_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF0000707F)) 
    \main_float64_addexit_0i_reg[63]_inv_i_2 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I1(\main_inst/main_101_102_reg_reg_n_0_[63] ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_10_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_11_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_20 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFAAAE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_21 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_23_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000004000000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_22 
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_23 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_24 
       (.I0(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFFE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_3 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_float64_addexit_0i13_out ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_15_n_0 ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_17_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_18_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    \main_float64_addexit_0i_reg[63]_inv_i_4 
       (.I0(\main_float64_addexit_0i_reg[62]_i_4_n_0 ),
        .I1(\main_inst/main_float64_addexit_0i121_out ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \main_float64_addexit_0i_reg[63]_inv_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \main_float64_addexit_0i_reg[63]_inv_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(main_158_160_reg),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \main_float64_addexit_0i_reg[63]_inv_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_20_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000020000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_8 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\roundAndPackFloat64_return_val_reg[63]_i_5_n_0 ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000001010100000)) 
    \main_float64_addexit_0i_reg[63]_inv_i_9 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_158_160_reg[62]_i_4_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[6]_i_1 
       (.I0(\main_float64_addexit_0i_reg[6]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[6]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[6]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[6]_i_2 
       (.I0(\main_float64_addexit_0i_reg[6]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [15]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[6]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[6] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [15]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[6]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[6]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [15]),
        .O(\main_float64_addexit_0i_reg[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[6]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[6] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [15]),
        .O(\main_float64_addexit_0i_reg[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[6]_i_6 
       (.I0(\main_inst/main_15_17 [15]),
        .I1(\main_inst/data5 [6]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[7]_i_1 
       (.I0(\main_float64_addexit_0i_reg[7]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[7]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[7]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[7]_i_10 
       (.I0(\main_inst/main_15_19_reg [14]),
        .I1(\main_inst/main_91_92 [14]),
        .O(\main_float64_addexit_0i_reg[7]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[7]_i_11 
       (.I0(\main_inst/main_15_19_reg [13]),
        .I1(\main_inst/main_91_92 [13]),
        .O(\main_float64_addexit_0i_reg[7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[7]_i_2 
       (.I0(\main_float64_addexit_0i_reg[7]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [16]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[7]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[7] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [16]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[7]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[7]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [16]),
        .O(\main_float64_addexit_0i_reg[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[7]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[7] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [16]),
        .O(\main_float64_addexit_0i_reg[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[7]_i_6 
       (.I0(\main_inst/main_15_17 [16]),
        .I1(\main_inst/data5 [7]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[7]_i_8 
       (.I0(\main_inst/main_15_19_reg [16]),
        .I1(\main_inst/main_91_92 [16]),
        .O(\main_float64_addexit_0i_reg[7]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_0i_reg[7]_i_9 
       (.I0(\main_inst/main_15_19_reg [15]),
        .I1(\main_inst/main_91_92 [15]),
        .O(\main_float64_addexit_0i_reg[7]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[8]_i_1 
       (.I0(\main_float64_addexit_0i_reg[8]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[8]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[8]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[8]_i_2 
       (.I0(\main_float64_addexit_0i_reg[8]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [17]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[8]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[8] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [17]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[8]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[8]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [17]),
        .O(\main_float64_addexit_0i_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[8]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[8] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [17]),
        .O(\main_float64_addexit_0i_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[8]_i_6 
       (.I0(\main_inst/main_15_17 [17]),
        .I1(\main_inst/data5 [8]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT4 #(
    .INIT(16'hFE0E)) 
    \main_float64_addexit_0i_reg[9]_i_1 
       (.I0(\main_float64_addexit_0i_reg[9]_i_2_n_0 ),
        .I1(\main_float64_addexit_0i_reg[9]_i_3_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_12_n_0 ),
        .I3(\main_float64_addexit_0i_reg[9]_i_4_n_0 ),
        .O(\main_float64_addexit_0i_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0300000022222222)) 
    \main_float64_addexit_0i_reg[9]_i_2 
       (.I0(\main_float64_addexit_0i_reg[9]_i_5_n_0 ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .I2(\main_float64_addexit_0i_reg[63]_inv_i_16_n_0 ),
        .I3(\main_inst/main_15_17 [18]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_22_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_21_n_0 ),
        .O(\main_float64_addexit_0i_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFBF8F8F800000000)) 
    \main_float64_addexit_0i_reg[9]_i_3 
       (.I0(\main_inst/main_101_102_reg_reg_n_0_[9] ),
        .I1(\main_float64_addexit_0i_reg[63]_inv_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_10_n_0 ),
        .I3(\main_inst/main_15_17 [18]),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_6_n_0 ),
        .I5(\main_float64_addexit_0i_reg[63]_inv_i_9_n_0 ),
        .O(\main_float64_addexit_0i_reg[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFDA800005500)) 
    \main_float64_addexit_0i_reg[9]_i_4 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_24_n_0 ),
        .I1(\main_float64_addexit_0i_reg[62]_i_5_n_0 ),
        .I2(\main_float64_addexit_0i_reg[62]_i_3_n_0 ),
        .I3(\main_float64_addexit_0i_reg[9]_i_6_n_0 ),
        .I4(\main_inst/main_float64_addexit_0i129_out ),
        .I5(\main_inst/main_15_17 [18]),
        .O(\main_float64_addexit_0i_reg[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE04)) 
    \main_float64_addexit_0i_reg[9]_i_5 
       (.I0(\main_float64_addexit_0i_reg[63]_inv_i_13_n_0 ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[9] ),
        .I2(\main_inst/main_float64_addexit_0i13_out ),
        .I3(\main_inst/main_15_17 [18]),
        .O(\main_float64_addexit_0i_reg[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hAAAAACA0)) 
    \main_float64_addexit_0i_reg[9]_i_6 
       (.I0(\main_inst/main_15_17 [18]),
        .I1(\main_inst/data5 [9]),
        .I2(\main_inst/main_float64_addexit_0i121_out ),
        .I3(\main_float64_addexit_0i_reg[63]_inv_i_8_n_0 ),
        .I4(\main_float64_addexit_0i_reg[63]_inv_i_7_n_0 ),
        .O(\main_float64_addexit_0i_reg[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[11]_i_7 
       (.CI(\main_float64_addexit_0i_reg_reg[7]_i_7_n_0 ),
        .CO(main_float64_addexit_0i_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [20:17]),
        .O(\main_inst/data5 [11:8]),
        .S({\main_float64_addexit_0i_reg[11]_i_8_n_0 ,\main_float64_addexit_0i_reg[11]_i_9_n_0 ,\main_float64_addexit_0i_reg[11]_i_10_n_0 ,\main_float64_addexit_0i_reg[11]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[15]_i_7 
       (.CI(main_float64_addexit_0i_reg_reg[3]),
        .CO({\main_float64_addexit_0i_reg_reg[15]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[15]_i_7_n_1 ,\main_float64_addexit_0i_reg_reg[15]_i_7_n_2 ,\main_float64_addexit_0i_reg_reg[15]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [24:21]),
        .O(\main_inst/data5 [15:12]),
        .S({\main_float64_addexit_0i_reg[15]_i_8_n_0 ,\main_float64_addexit_0i_reg[15]_i_9_n_0 ,\main_float64_addexit_0i_reg[15]_i_10_n_0 ,\main_float64_addexit_0i_reg[15]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[19]_i_7 
       (.CI(\main_float64_addexit_0i_reg_reg[15]_i_7_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[19]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[19]_i_7_n_1 ,\main_float64_addexit_0i_reg_reg[19]_i_7_n_2 ,\main_float64_addexit_0i_reg_reg[19]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [28:25]),
        .O(\main_inst/data5 [19:16]),
        .S({\main_float64_addexit_0i_reg[19]_i_8_n_0 ,\main_float64_addexit_0i_reg[19]_i_9_n_0 ,\main_float64_addexit_0i_reg[19]_i_10_n_0 ,\main_float64_addexit_0i_reg[19]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[23]_i_7 
       (.CI(\main_float64_addexit_0i_reg_reg[19]_i_7_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[23]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[23]_i_7_n_1 ,\main_float64_addexit_0i_reg_reg[23]_i_7_n_2 ,\main_float64_addexit_0i_reg_reg[23]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [32:29]),
        .O(\main_inst/data5 [23:20]),
        .S({\main_float64_addexit_0i_reg[23]_i_8_n_0 ,\main_float64_addexit_0i_reg[23]_i_9_n_0 ,\main_float64_addexit_0i_reg[23]_i_10_n_0 ,\main_float64_addexit_0i_reg[23]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[32]_i_5 
       (.CI(\main_float64_addexit_0i_reg_reg[32]_i_6_n_0 ),
        .CO({\main_inst/data5 [32],\main_float64_addexit_0i_reg_reg[32]_i_5_n_1 ,\main_float64_addexit_0i_reg_reg[32]_i_5_n_2 ,\main_float64_addexit_0i_reg_reg[32]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [40:37]),
        .O(\main_inst/data5 [31:28]),
        .S({\main_float64_addexit_0i_reg[32]_i_7_n_0 ,\main_float64_addexit_0i_reg[32]_i_8_n_0 ,\main_float64_addexit_0i_reg[32]_i_9_n_0 ,\main_float64_addexit_0i_reg[32]_i_10_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[32]_i_6 
       (.CI(\main_float64_addexit_0i_reg_reg[23]_i_7_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[32]_i_6_n_0 ,\main_float64_addexit_0i_reg_reg[32]_i_6_n_1 ,\main_float64_addexit_0i_reg_reg[32]_i_6_n_2 ,\main_float64_addexit_0i_reg_reg[32]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [36:33]),
        .O(\main_inst/data5 [27:24]),
        .S({\main_float64_addexit_0i_reg[32]_i_11_n_0 ,\main_float64_addexit_0i_reg[32]_i_12_n_0 ,\main_float64_addexit_0i_reg[32]_i_13_n_0 ,\main_float64_addexit_0i_reg[32]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[3]_i_7 
       (.CI(\<const0>__0__0 ),
        .CO({\main_float64_addexit_0i_reg_reg[3]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[3]_i_7_n_1 ,\main_float64_addexit_0i_reg_reg[3]_i_7_n_2 ,\main_float64_addexit_0i_reg_reg[3]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [12:9]),
        .O({\main_inst/data5 [3:1],\main_float64_addexit_0i_reg_reg[3]_i_7_n_7 }),
        .S({\main_float64_addexit_0i_reg[3]_i_8_n_0 ,\main_float64_addexit_0i_reg[3]_i_9_n_0 ,\main_float64_addexit_0i_reg[3]_i_10_n_0 ,\main_inst/data5 [0]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[62]_i_11 
       (.CI(\main_float64_addexit_0i_reg_reg[62]_i_12_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[62]_i_11_n_0 ,\main_float64_addexit_0i_reg_reg[62]_i_11_n_1 ,\main_float64_addexit_0i_reg_reg[62]_i_11_n_2 ,\main_float64_addexit_0i_reg_reg[62]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[62]_i_12 
       (.CI(\main_float64_addexit_0i_reg_reg[62]_i_13_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[62]_i_12_n_0 ,\main_float64_addexit_0i_reg_reg[62]_i_12_n_1 ,\main_float64_addexit_0i_reg_reg[62]_i_12_n_2 ,\main_float64_addexit_0i_reg_reg[62]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const1>__0__0 ,\main_float64_addexit_0i_reg[62]_i_14_n_0 ,\main_float64_addexit_0i_reg[62]_i_15_n_0 ,\main_float64_addexit_0i_reg[62]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[62]_i_13 
       (.CI(\main_float64_addexit_0i_reg_reg[62]_i_17_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[62]_i_13_n_0 ,\main_float64_addexit_0i_reg_reg[62]_i_13_n_1 ,\main_float64_addexit_0i_reg_reg[62]_i_13_n_2 ,\main_float64_addexit_0i_reg_reg[62]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_0i_reg[62]_i_18_n_0 ,\main_float64_addexit_0i_reg[62]_i_19_n_0 ,\main_float64_addexit_0i_reg[62]_i_20_n_0 ,\main_float64_addexit_0i_reg[62]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[62]_i_17 
       (.CI(\<const0>__0__0 ),
        .CO({\main_float64_addexit_0i_reg_reg[62]_i_17_n_0 ,\main_float64_addexit_0i_reg_reg[62]_i_17_n_1 ,\main_float64_addexit_0i_reg_reg[62]_i_17_n_2 ,\main_float64_addexit_0i_reg_reg[62]_i_17_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_0i_reg[62]_i_22_n_0 ,\main_float64_addexit_0i_reg[62]_i_23_n_0 ,\main_float64_addexit_0i_reg[62]_i_24_n_0 ,\main_float64_addexit_0i_reg[62]_i_25_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[62]_i_7 
       (.CI(\main_float64_addexit_0i_reg_reg[62]_i_11_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[62]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[62]_i_7_n_1 ,\main_inst/main_23_24 ,\main_float64_addexit_0i_reg_reg[62]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_0i_reg_reg[7]_i_7 
       (.CI(\main_float64_addexit_0i_reg_reg[3]_i_7_n_0 ),
        .CO({\main_float64_addexit_0i_reg_reg[7]_i_7_n_0 ,\main_float64_addexit_0i_reg_reg[7]_i_7_n_1 ,\main_float64_addexit_0i_reg_reg[7]_i_7_n_2 ,\main_float64_addexit_0i_reg_reg[7]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/main_15_19_reg [16:13]),
        .O(\main_inst/data5 [7:4]),
        .S({\main_float64_addexit_0i_reg[7]_i_8_n_0 ,\main_float64_addexit_0i_reg[7]_i_9_n_0 ,\main_float64_addexit_0i_reg[7]_i_10_n_0 ,\main_float64_addexit_0i_reg[7]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004000000000000)) 
    \main_float64_addexit_218_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\return_val[31]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_inst/main_float64_addexit_218_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_10 
       (.I0(\main_inst/main_float64_addexit_0i_reg [57]),
        .I1(\main_inst/main_float64_addexit_0i_reg [59]),
        .I2(\main_inst/main_float64_addexit_0i_reg [58]),
        .O(main_float64_addexit_218_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_11 
       (.I0(\main_inst/main_float64_addexit_0i_reg [54]),
        .I1(\main_inst/main_float64_addexit_0i_reg [56]),
        .I2(\main_inst/main_float64_addexit_0i_reg [55]),
        .O(\main_float64_addexit_218_reg[3]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_12 
       (.I0(\main_inst/main_float64_addexit_0i_reg [51]),
        .I1(\main_inst/main_float64_addexit_0i_reg [53]),
        .I2(\main_inst/main_float64_addexit_0i_reg [52]),
        .O(\main_float64_addexit_218_reg[3]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_13 
       (.I0(\main_inst/main_float64_addexit_0i_reg [48]),
        .I1(\main_inst/main_float64_addexit_0i_reg [50]),
        .I2(\main_inst/main_float64_addexit_0i_reg [49]),
        .O(\main_float64_addexit_218_reg[3]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_15 
       (.I0(\main_inst/main_float64_addexit_0i_reg [45]),
        .I1(\main_inst/main_float64_addexit_0i_reg [47]),
        .I2(\main_inst/main_float64_addexit_0i_reg [46]),
        .O(\main_float64_addexit_218_reg[3]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_16 
       (.I0(\main_inst/main_float64_addexit_0i_reg [42]),
        .I1(\main_inst/main_float64_addexit_0i_reg [44]),
        .I2(\main_inst/main_float64_addexit_0i_reg [43]),
        .O(\main_float64_addexit_218_reg[3]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_17 
       (.I0(\main_inst/main_float64_addexit_0i_reg [39]),
        .I1(\main_inst/main_float64_addexit_0i_reg [41]),
        .I2(\main_inst/main_float64_addexit_0i_reg [40]),
        .O(\main_float64_addexit_218_reg[3]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_18 
       (.I0(\main_inst/main_float64_addexit_0i_reg [36]),
        .I1(\main_inst/main_float64_addexit_0i_reg [38]),
        .I2(\main_inst/main_float64_addexit_0i_reg [37]),
        .O(\main_float64_addexit_218_reg[3]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_20 
       (.I0(\main_inst/main_float64_addexit_0i_reg [33]),
        .I1(\main_inst/main_float64_addexit_0i_reg [35]),
        .I2(\main_inst/main_float64_addexit_0i_reg [34]),
        .O(\main_float64_addexit_218_reg[3]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h09000009)) 
    \main_float64_addexit_218_reg[3]_i_21 
       (.I0(\main_inst/main_float64_addexit_0i_reg [30]),
        .I1(memory_controller_out_a[30]),
        .I2(\main_inst/main_float64_addexit_0i_reg [32]),
        .I3(memory_controller_out_a[31]),
        .I4(\main_inst/main_float64_addexit_0i_reg [31]),
        .O(\main_float64_addexit_218_reg[3]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_22 
       (.I0(\main_inst/main_float64_addexit_0i_reg [27]),
        .I1(memory_controller_out_a[27]),
        .I2(memory_controller_out_a[29]),
        .I3(\main_inst/main_float64_addexit_0i_reg [29]),
        .I4(memory_controller_out_a[28]),
        .I5(\main_inst/main_float64_addexit_0i_reg [28]),
        .O(\main_float64_addexit_218_reg[3]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_23 
       (.I0(\main_inst/main_float64_addexit_0i_reg [24]),
        .I1(memory_controller_out_a[24]),
        .I2(memory_controller_out_a[26]),
        .I3(\main_inst/main_float64_addexit_0i_reg [26]),
        .I4(memory_controller_out_a[25]),
        .I5(\main_inst/main_float64_addexit_0i_reg [25]),
        .O(\main_float64_addexit_218_reg[3]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_25 
       (.I0(\main_inst/main_float64_addexit_0i_reg [21]),
        .I1(memory_controller_out_a[21]),
        .I2(memory_controller_out_a[23]),
        .I3(\main_inst/main_float64_addexit_0i_reg [23]),
        .I4(memory_controller_out_a[22]),
        .I5(\main_inst/main_float64_addexit_0i_reg [22]),
        .O(\main_float64_addexit_218_reg[3]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_26 
       (.I0(\main_inst/main_float64_addexit_0i_reg [18]),
        .I1(memory_controller_out_a[18]),
        .I2(memory_controller_out_a[20]),
        .I3(\main_inst/main_float64_addexit_0i_reg [20]),
        .I4(memory_controller_out_a[19]),
        .I5(\main_inst/main_float64_addexit_0i_reg [19]),
        .O(\main_float64_addexit_218_reg[3]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_27 
       (.I0(\main_inst/main_float64_addexit_0i_reg [15]),
        .I1(memory_controller_out_a[15]),
        .I2(memory_controller_out_a[17]),
        .I3(\main_inst/main_float64_addexit_0i_reg [17]),
        .I4(memory_controller_out_a[16]),
        .I5(\main_inst/main_float64_addexit_0i_reg [16]),
        .O(\main_float64_addexit_218_reg[3]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_28 
       (.I0(\main_inst/main_float64_addexit_0i_reg [12]),
        .I1(memory_controller_out_a[12]),
        .I2(memory_controller_out_a[14]),
        .I3(\main_inst/main_float64_addexit_0i_reg [14]),
        .I4(memory_controller_out_a[13]),
        .I5(\main_inst/main_float64_addexit_0i_reg [13]),
        .O(\main_float64_addexit_218_reg[3]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_29 
       (.I0(\main_inst/main_float64_addexit_0i_reg [9]),
        .I1(memory_controller_out_a[9]),
        .I2(memory_controller_out_a[11]),
        .I3(\main_inst/main_float64_addexit_0i_reg [11]),
        .I4(memory_controller_out_a[10]),
        .I5(\main_inst/main_float64_addexit_0i_reg [10]),
        .O(\main_float64_addexit_218_reg[3]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_30 
       (.I0(\main_inst/main_float64_addexit_0i_reg [6]),
        .I1(memory_controller_out_a[6]),
        .I2(memory_controller_out_a[8]),
        .I3(\main_inst/main_float64_addexit_0i_reg [8]),
        .I4(memory_controller_out_a[7]),
        .I5(\main_inst/main_float64_addexit_0i_reg [7]),
        .O(\main_float64_addexit_218_reg[3]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_31 
       (.I0(\main_inst/main_float64_addexit_0i_reg [3]),
        .I1(memory_controller_out_a[3]),
        .I2(memory_controller_out_a[5]),
        .I3(\main_inst/main_float64_addexit_0i_reg [5]),
        .I4(memory_controller_out_a[4]),
        .I5(\main_inst/main_float64_addexit_0i_reg [4]),
        .O(\main_float64_addexit_218_reg[3]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9009000000009009)) 
    \main_float64_addexit_218_reg[3]_i_32 
       (.I0(\main_inst/main_float64_addexit_0i_reg [0]),
        .I1(memory_controller_out_a[0]),
        .I2(memory_controller_out_a[2]),
        .I3(\main_inst/main_float64_addexit_0i_reg [2]),
        .I4(memory_controller_out_a[1]),
        .I5(\main_inst/main_float64_addexit_0i_reg [1]),
        .O(\main_float64_addexit_218_reg[3]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_float64_addexit_218_reg[3]_i_6 
       (.I0(\main_inst/CI ),
        .I1(\main_inst/main_1_main_result02_reg_reg [0]),
        .O(\main_float64_addexit_218_reg[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_float64_addexit_218_reg[3]_i_8 
       (.I0(\main_inst/main_float64_addexit_0i_reg [60]),
        .I1(\main_inst/main_float64_addexit_0i_reg [62]),
        .I2(\main_inst/main_float64_addexit_0i_reg [61]),
        .O(\main_float64_addexit_218_reg[3]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[11]_i_1 
       (.CI(\main_float64_addexit_218_reg_reg[7]_i_1_n_0 ),
        .CO(main_float64_addexit_218_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [11:8]),
        .S(\main_inst/main_1_main_result02_reg_reg [11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[15]_i_1 
       (.CI(main_float64_addexit_218_reg_reg[3]),
        .CO({\main_float64_addexit_218_reg_reg[15]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[15]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[15]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [15:12]),
        .S(\main_inst/main_1_main_result02_reg_reg [15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[19]_i_1 
       (.CI(\main_float64_addexit_218_reg_reg[15]_i_1_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[19]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[19]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[19]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [19:16]),
        .S(\main_inst/main_1_main_result02_reg_reg [19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[23]_i_1 
       (.CI(\main_float64_addexit_218_reg_reg[19]_i_1_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[23]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[23]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[23]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [23:20]),
        .S(\main_inst/main_1_main_result02_reg_reg [23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[27]_i_1 
       (.CI(\main_float64_addexit_218_reg_reg[23]_i_1_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[27]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[27]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[27]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [27:24]),
        .S(\main_inst/main_1_main_result02_reg_reg [27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[31]_i_2 
       (.CI(\main_float64_addexit_218_reg_reg[27]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [31:28]),
        .S(\main_inst/main_1_main_result02_reg_reg [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/CI }),
        .O(\main_inst/main_float64_addexit_218 [3:0]),
        .S({\main_inst/main_1_main_result02_reg_reg [3:1],\main_float64_addexit_218_reg[3]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_14 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_19_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_14_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_14_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_14_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_14_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_218_reg[3]_i_20_n_0 ,\main_float64_addexit_218_reg[3]_i_21_n_0 ,\main_float64_addexit_218_reg[3]_i_22_n_0 ,\main_float64_addexit_218_reg[3]_i_23_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_19 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_24_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_19_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_19_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_19_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_218_reg[3]_i_25_n_0 ,\main_float64_addexit_218_reg[3]_i_26_n_0 ,\main_float64_addexit_218_reg[3]_i_27_n_0 ,\main_float64_addexit_218_reg[3]_i_28_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_2 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_7_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_2_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_2_n_1 ,\main_inst/CI ,\main_float64_addexit_218_reg_reg[3]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_float64_addexit_0i_reg_reg ,\main_float64_addexit_218_reg[3]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_24 
       (.CI(\<const0>__0__0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_24_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_24_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_24_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_24_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_218_reg[3]_i_29_n_0 ,\main_float64_addexit_218_reg[3]_i_30_n_0 ,\main_float64_addexit_218_reg[3]_i_31_n_0 ,\main_float64_addexit_218_reg[3]_i_32_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_7 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_9_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_7_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_7_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_7_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({main_float64_addexit_218_reg,\main_float64_addexit_218_reg[3]_i_11_n_0 ,\main_float64_addexit_218_reg[3]_i_12_n_0 ,\main_float64_addexit_218_reg[3]_i_13_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[3]_i_9 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_14_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[3]_i_9_n_0 ,\main_float64_addexit_218_reg_reg[3]_i_9_n_1 ,\main_float64_addexit_218_reg_reg[3]_i_9_n_2 ,\main_float64_addexit_218_reg_reg[3]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .S({\main_float64_addexit_218_reg[3]_i_15_n_0 ,\main_float64_addexit_218_reg[3]_i_16_n_0 ,\main_float64_addexit_218_reg[3]_i_17_n_0 ,\main_float64_addexit_218_reg[3]_i_18_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_218_reg_reg[7]_i_1 
       (.CI(\main_float64_addexit_218_reg_reg[3]_i_1_n_0 ),
        .CO({\main_float64_addexit_218_reg_reg[7]_i_1_n_0 ,\main_float64_addexit_218_reg_reg[7]_i_1_n_1 ,\main_float64_addexit_218_reg_reg[7]_i_1_n_2 ,\main_float64_addexit_218_reg_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_218 [7:4]),
        .S(\main_inst/main_1_main_result02_reg_reg [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \main_float64_addexit_220_reg[0]_i_1 
       (.I0(\main_inst/main_1_scevgep_reg1 [3]),
        .O(\main_inst/main_float64_addexit_220 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \main_float64_addexit_220_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(main_float64_addexit_220_reg),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/main_float64_addexit_220_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \main_float64_addexit_220_reg[31]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .O(main_float64_addexit_220_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[12]_i_1 
       (.CI(\main_float64_addexit_220_reg_reg[8]_i_1_n_0 ),
        .CO(main_float64_addexit_220_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [12:9]),
        .S(\main_inst/main_1_scevgep_reg1 [15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[16]_i_1 
       (.CI(main_float64_addexit_220_reg_reg[3]),
        .CO({\main_float64_addexit_220_reg_reg[16]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[16]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[16]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[16]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [16:13]),
        .S(\main_inst/main_1_scevgep_reg1 [19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[20]_i_1 
       (.CI(\main_float64_addexit_220_reg_reg[16]_i_1_n_0 ),
        .CO({\main_float64_addexit_220_reg_reg[20]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[20]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[20]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[20]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [20:17]),
        .S(\main_inst/main_1_scevgep_reg1 [23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[24]_i_1 
       (.CI(\main_float64_addexit_220_reg_reg[20]_i_1_n_0 ),
        .CO({\main_float64_addexit_220_reg_reg[24]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[24]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[24]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[24]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [24:21]),
        .S(\main_inst/main_1_scevgep_reg1 [27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[28]_i_1 
       (.CI(\main_float64_addexit_220_reg_reg[24]_i_1_n_0 ),
        .CO({\main_float64_addexit_220_reg_reg[28]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[28]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[28]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[28]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [28:25]),
        .S(\main_inst/main_1_scevgep_reg1 [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[31]_i_2 
       (.CI(\main_float64_addexit_220_reg_reg[28]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_float64_addexit_220_reg_reg[31]_i_2_n_4 ,\main_inst/main_float64_addexit_220 [31:29]}),
        .S({\<const0>__0__0 ,\main_inst/main_1_2_reg_reg_n_0_[31] ,\main_inst/main_1_2_reg_reg_n_0_[30] ,\main_inst/main_1_2_reg_reg_n_0_ }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[4]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\main_float64_addexit_220_reg_reg[4]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[4]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[4]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[4]_i_1_n_3 }),
        .CYINIT(\main_inst/main_1_scevgep_reg1 [3]),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [4:1]),
        .S(\main_inst/main_1_scevgep_reg1 [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_float64_addexit_220_reg_reg[8]_i_1 
       (.CI(\main_float64_addexit_220_reg_reg[4]_i_1_n_0 ),
        .CO({\main_float64_addexit_220_reg_reg[8]_i_1_n_0 ,\main_float64_addexit_220_reg_reg[8]_i_1_n_1 ,\main_float64_addexit_220_reg_reg[8]_i_1_n_2 ,\main_float64_addexit_220_reg_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_float64_addexit_220 [8:5]),
        .S(\main_inst/main_1_scevgep_reg1 [11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h4000)) 
    main_float64_addexit_exitcond1_reg_i_1
       (.I0(main_float64_addexit_exitcond1_reg_i_2_n_0),
        .I1(main_float64_addexit_exitcond1_reg_i_3_n_0),
        .I2(main_float64_addexit_exitcond1_reg_i_4_n_0),
        .I3(main_float64_addexit_exitcond1_reg_i_5_n_0),
        .O(\main_inst/main_float64_addexit_exitcond1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFEFFFF)) 
    main_float64_addexit_exitcond1_reg_i_2
       (.I0(\main_inst/main_float64_addexit_220 [16]),
        .I1(\main_inst/main_float64_addexit_220 [17]),
        .I2(\main_inst/main_float64_addexit_220 [18]),
        .I3(\main_inst/main_float64_addexit_220 [19]),
        .I4(main_float64_addexit_exitcond1_reg_i_6_n_0),
        .O(main_float64_addexit_exitcond1_reg_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    main_float64_addexit_exitcond1_reg_i_3
       (.I0(\main_inst/main_float64_addexit_220 [28]),
        .I1(\main_inst/main_float64_addexit_220 [29]),
        .I2(\main_inst/main_float64_addexit_220 [31]),
        .I3(\main_inst/main_float64_addexit_220 [30]),
        .I4(main_float64_addexit_exitcond1_reg_i_7_n_0),
        .O(main_float64_addexit_exitcond1_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    main_float64_addexit_exitcond1_reg_i_4
       (.I0(\main_inst/main_float64_addexit_220 [12]),
        .I1(\main_inst/main_float64_addexit_220 [13]),
        .I2(\main_inst/main_float64_addexit_220 [14]),
        .I3(\main_inst/main_float64_addexit_220 [15]),
        .I4(main_float64_addexit_exitcond1_reg_i_8_n_0),
        .O(main_float64_addexit_exitcond1_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000004)) 
    main_float64_addexit_exitcond1_reg_i_5
       (.I0(\main_inst/main_float64_addexit_220 [4]),
        .I1(\main_inst/main_1_scevgep_reg1 [3]),
        .I2(\main_inst/main_float64_addexit_220 [6]),
        .I3(\main_inst/main_float64_addexit_220 [7]),
        .I4(main_float64_addexit_exitcond1_reg_i_9_n_0),
        .O(main_float64_addexit_exitcond1_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0001)) 
    main_float64_addexit_exitcond1_reg_i_6
       (.I0(\main_inst/main_float64_addexit_220 [23]),
        .I1(\main_inst/main_float64_addexit_220 [22]),
        .I2(\main_inst/main_float64_addexit_220 [21]),
        .I3(\main_inst/main_float64_addexit_220 [20]),
        .O(main_float64_addexit_exitcond1_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    main_float64_addexit_exitcond1_reg_i_7
       (.I0(\main_inst/main_float64_addexit_220 [25]),
        .I1(\main_inst/main_float64_addexit_220 [24]),
        .I2(\main_inst/main_float64_addexit_220 [27]),
        .I3(\main_inst/main_float64_addexit_220 [26]),
        .O(main_float64_addexit_exitcond1_reg_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFFE)) 
    main_float64_addexit_exitcond1_reg_i_8
       (.I0(\main_inst/main_float64_addexit_220 [9]),
        .I1(\main_inst/main_float64_addexit_220 [8]),
        .I2(\main_inst/main_float64_addexit_220 [11]),
        .I3(\main_inst/main_float64_addexit_220 [10]),
        .O(main_float64_addexit_exitcond1_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    main_float64_addexit_exitcond1_reg_i_9
       (.I0(\main_inst/main_float64_addexit_220 [2]),
        .I1(\main_inst/main_float64_addexit_220 [1]),
        .I2(\main_inst/main_float64_addexit_220 [5]),
        .I3(\main_inst/main_float64_addexit_220 [3]),
        .O(main_float64_addexit_exitcond1_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[0] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [0]),
        .Q(\main_inst/cur_state_reg_n_0_ ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "cur_state_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[1] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [1]),
        .Q(\main_inst/cur_state_reg_n_0_[1] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "cur_state_reg[1]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[1]_rep 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\cur_state[1]_rep_i_1_n_0 ),
        .Q(\main_inst/cur_state_reg ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[2] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [2]),
        .Q(\main_inst/cur_state_reg_n_0_[2] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[3] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [3]),
        .Q(\main_inst/cur_state_reg_n_0_[3] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[4] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [4]),
        .Q(\main_inst/cur_state_reg_n_0_[4] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[5] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\cur_state[5]_i_1_n_0 ),
        .Q(\main_inst/cur_state_reg_n_0_[5] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "cur_state_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[6] 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [6]),
        .Q(\main_inst/cur_state_reg_n_0_[6] ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* ORIG_CELL_NAME = "cur_state_reg[6]" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/cur_state_reg[6]_rep 
       (.C(clk),
        .CE(\main_inst/cur_state ),
        .D(\main_inst/next_state [6]),
        .Q(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAAAAC)) 
    \main_inst/finish_i_1 
       (.I0(\main_inst/roundAndPackFloat64_finish ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\main_inst/finish_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/finish_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(finish_i_1_n_0),
        .Q(finish),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [0]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [10]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [11]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [12]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [13]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [14]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [15]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [16]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [17]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [18]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [19]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [1]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [20]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [21]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [22]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [23]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [24]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [25]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [26]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [27]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [28]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [29]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [2]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [30]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [31]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [32]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [33]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [34]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [35]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [36]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [37]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [38]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [39]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [3]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [40]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [41]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [42]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [43]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [44]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [45]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [46]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [47]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [48]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [49]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [4]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [50]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [51]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [52]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [53]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [54]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [55]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [56]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [57]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [58]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [59]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [5]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [60]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [61]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [62]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [63]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [6]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [7]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [8]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_102_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_101_102_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [9]),
        .Q(\main_inst/main_101_102_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[3]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[11]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[11]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[15]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[15]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[15]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[15]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[19]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[19]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[19]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[19]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[3]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[23]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[23]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[23]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[23]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[27]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[27]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[27]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[27]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[31]_i_2_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[31]_i_2_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[3]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[31]_i_2_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[31]_i_2_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[3]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[7]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[7]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[7]_i_1_n_5 ),
        .Q(\main_inst/main_101_zExp1ii_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[7]_i_1_n_4 ),
        .Q(\main_inst/main_101_zExp1ii_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[11]_i_1_n_7 ),
        .Q(\main_inst/main_101_zExp1ii_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zExp1ii_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zExp1ii_reg_reg[11]_i_1_n_6 ),
        .Q(\main_inst/main_101_zExp1ii_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[12]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[12]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[12]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[16]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[16]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[16]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[16]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[20]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[20]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[20]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [1]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[1] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[20]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[24]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[24]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[24]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[24]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[28]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[28]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[28]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[28]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[32]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [2]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[2] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[32]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[32]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[32]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[36]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[36]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[36]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[36]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[40]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[40]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[40]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [3]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[3] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[40]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[44]_i_1_n_7 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[44]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[44]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[44]_i_1_n_4 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [4]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[4] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [5]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[5] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[63]_i_1_n_6 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg_reg[63]_i_1_n_5 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [6]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[6] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [7]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[7] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_ii_reg [8]),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[8] ),
        .R(\main_101_zSig0i12i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_101_zSig0i12i_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_101_zSig0i12i_reg ),
        .D(\main_101_zSig0i12i_reg[9]_i_1_n_0 ),
        .Q(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [9]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [10]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [11]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [12]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [13]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [14]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [15]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [16]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [17]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [18]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [19]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [20]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [21]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [22]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [23]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [24]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [25]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [26]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [27]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [28]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [29]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [30]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [31]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [32]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [33]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [34]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [35]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [36]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [37]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [38]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [39]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_105_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_15_17 [40]),
        .Q(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [10]),
        .Q(\main_inst/main_103_107_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [11]),
        .Q(\main_inst/main_103_107_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [12]),
        .Q(\main_inst/main_103_107_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [13]),
        .Q(\main_inst/main_103_107_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [14]),
        .Q(\main_inst/main_103_107_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [15]),
        .Q(\main_inst/main_103_107_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [16]),
        .Q(\main_inst/main_103_107_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [17]),
        .Q(\main_inst/main_103_107_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [18]),
        .Q(\main_inst/main_103_107_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [19]),
        .Q(\main_inst/main_103_107_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [20]),
        .Q(\main_inst/main_103_107_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [21]),
        .Q(\main_inst/main_103_107_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [22]),
        .Q(\main_inst/main_103_107_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [23]),
        .Q(\main_inst/main_103_107_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [24]),
        .Q(\main_inst/main_103_107_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [25]),
        .Q(\main_inst/main_103_107_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [26]),
        .Q(\main_inst/main_103_107_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [27]),
        .Q(\main_inst/main_103_107_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [28]),
        .Q(\main_inst/main_103_107_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [29]),
        .Q(\main_inst/main_103_107_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [30]),
        .Q(\main_inst/main_103_107_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [31]),
        .Q(\main_inst/main_103_107_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [32]),
        .Q(\main_inst/main_103_107_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [33]),
        .Q(\main_inst/main_103_107_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [34]),
        .Q(\main_inst/main_103_107_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [35]),
        .Q(\main_inst/main_103_107_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [36]),
        .Q(\main_inst/main_103_107_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [37]),
        .Q(\main_inst/main_103_107_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [38]),
        .Q(\main_inst/main_103_107_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [39]),
        .Q(\main_inst/main_103_107_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [40]),
        .Q(\main_inst/main_103_107_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_103_107_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_103_105_reg ),
        .D(\main_inst/main_103_107 [41]),
        .Q(\main_inst/main_103_107_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_121_aExp0ii_reg_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(main_121_aExp0ii_reg),
        .Q(\main_inst/main_121_aExp0ii_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_121_bExp0ii_reg_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(main_121_bExp0ii_reg),
        .Q(\main_inst/main_121_bExp0ii_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_ ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_139_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .Q(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_141_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(ONE_10),
        .Q(\main_inst/main_136_141_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_141_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(ONE_8),
        .Q(\main_inst/main_136_141_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_141_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(ONE_7),
        .Q(\main_inst/main_136_141_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_141_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(ONE_12),
        .Q(\main_inst/main_136_141_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_141_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(ONE_11),
        .Q(\main_inst/main_136_141_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_136_expDiff0ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_136_139_reg ),
        .D(main_136_expDiff0ii_reg_reg),
        .Q(\main_inst/main_136_expDiff0ii_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(main_158_159_reg),
        .Q(\main_inst/main_158_159_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [10]),
        .Q(\main_inst/main_158_159_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [11]),
        .Q(\main_inst/main_158_159_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [12]),
        .Q(\main_inst/main_158_159_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [13]),
        .Q(\main_inst/main_158_159_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [14]),
        .Q(\main_inst/main_158_159_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [15]),
        .Q(\main_inst/main_158_159_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [16]),
        .Q(\main_inst/main_158_159_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [17]),
        .Q(\main_inst/main_158_159_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [18]),
        .Q(\main_inst/main_158_159_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [19]),
        .Q(\main_inst/main_158_159_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [20]),
        .Q(\main_inst/main_158_159_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [21]),
        .Q(\main_inst/main_158_159_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [22]),
        .Q(\main_inst/main_158_159_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [23]),
        .Q(\main_inst/main_158_159_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [24]),
        .Q(\main_inst/main_158_159_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [25]),
        .Q(\main_inst/main_158_159_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [26]),
        .Q(\main_inst/main_158_159_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [27]),
        .Q(\main_inst/main_158_159_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [28]),
        .Q(\main_inst/main_158_159_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [29]),
        .Q(\main_inst/main_158_159_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [30]),
        .Q(\main_inst/main_158_159_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [31]),
        .Q(\main_inst/main_158_159_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [32]),
        .Q(\main_inst/main_158_159_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [33]),
        .Q(\main_inst/main_158_159_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [34]),
        .Q(\main_inst/main_158_159_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [35]),
        .Q(\main_inst/main_158_159_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [36]),
        .Q(\main_inst/main_158_159_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [37]),
        .Q(\main_inst/main_158_159_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [38]),
        .Q(\main_inst/main_158_159_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [39]),
        .Q(\main_inst/main_158_159_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [40]),
        .Q(\main_inst/main_158_159_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_159 [41]),
        .Q(\main_inst/main_158_159_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_159_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_158_159_reg[9]_i_1_n_0 ),
        .Q(\main_inst/main_158_159_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [10]),
        .Q(\main_inst/main_158_160_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [11]),
        .Q(\main_inst/main_158_160_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [12]),
        .Q(\main_inst/main_158_160_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [13]),
        .Q(\main_inst/main_158_160_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [14]),
        .Q(\main_inst/main_158_160_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [15]),
        .Q(\main_inst/main_158_160_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [16]),
        .Q(\main_inst/main_158_160_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [17]),
        .Q(\main_inst/main_158_160_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [18]),
        .Q(\main_inst/main_158_160_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [19]),
        .Q(\main_inst/main_158_160_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [20]),
        .Q(\main_inst/main_158_160_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [21]),
        .Q(\main_inst/main_158_160_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [22]),
        .Q(\main_inst/main_158_160_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [23]),
        .Q(\main_inst/main_158_160_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [24]),
        .Q(\main_inst/main_158_160_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [25]),
        .Q(\main_inst/main_158_160_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [26]),
        .Q(\main_inst/main_158_160_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [27]),
        .Q(\main_inst/main_158_160_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [28]),
        .Q(\main_inst/main_158_160_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [29]),
        .Q(\main_inst/main_158_160_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [30]),
        .Q(\main_inst/main_158_160_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [31]),
        .Q(\main_inst/main_158_160_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [32]),
        .Q(\main_inst/main_158_160_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [33]),
        .Q(\main_inst/main_158_160_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [34]),
        .Q(\main_inst/main_158_160_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [35]),
        .Q(\main_inst/main_158_160_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [36]),
        .Q(\main_inst/main_158_160_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [37]),
        .Q(\main_inst/main_158_160_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [38]),
        .Q(\main_inst/main_158_160_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [39]),
        .Q(\main_inst/main_158_160_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [40]),
        .Q(\main_inst/main_158_160_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_103_107_reg [41]),
        .Q(\main_inst/main_158_160_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_160_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(\main_inst/main_158_160 ),
        .Q(\main_inst/main_158_160_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_158_bExp1ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_158_bExp1ii_reg ),
        .D(main_158_bExp1ii_reg),
        .Q(\main_inst/main_158_bExp1ii_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [10]),
        .Q(\main_inst/main_91_92 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [11]),
        .Q(\main_inst/main_91_92 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [12]),
        .Q(\main_inst/main_91_92 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [13]),
        .Q(\main_inst/main_91_92 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [14]),
        .Q(\main_inst/main_91_92 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [15]),
        .Q(\main_inst/main_91_92 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [16]),
        .Q(\main_inst/main_91_92 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [17]),
        .Q(\main_inst/main_91_92 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [18]),
        .Q(\main_inst/main_91_92 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [19]),
        .Q(\main_inst/main_91_92 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [20]),
        .Q(\main_inst/main_91_92 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [21]),
        .Q(\main_inst/main_91_92 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [22]),
        .Q(\main_inst/main_91_92 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [23]),
        .Q(\main_inst/main_91_92 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [24]),
        .Q(\main_inst/main_91_92 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [25]),
        .Q(\main_inst/main_91_92 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [26]),
        .Q(\main_inst/main_91_92 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [27]),
        .Q(\main_inst/main_91_92 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [28]),
        .Q(\main_inst/main_91_92 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [29]),
        .Q(\main_inst/main_91_92 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [30]),
        .Q(\main_inst/main_91_92 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [31]),
        .Q(\main_inst/main_91_92 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [32]),
        .Q(\main_inst/main_91_92 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [33]),
        .Q(\main_inst/main_91_92 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [34]),
        .Q(\main_inst/main_91_92 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [35]),
        .Q(\main_inst/main_91_92 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [36]),
        .Q(\main_inst/main_91_92 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [37]),
        .Q(\main_inst/main_91_92 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [38]),
        .Q(\main_inst/main_91_92 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [39]),
        .Q(\main_inst/main_91_92 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [40]),
        .Q(\main_inst/main_91_92 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_17_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_15_17 [9]),
        .Q(\main_inst/main_91_92 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [11]),
        .Q(\main_inst/main_15_19_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [12]),
        .Q(\main_inst/main_15_19_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [13]),
        .Q(\main_inst/main_15_19_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [14]),
        .Q(\main_inst/main_15_19_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [15]),
        .Q(\main_inst/main_15_19_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [16]),
        .Q(\main_inst/main_15_19_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [17]),
        .Q(\main_inst/main_15_19_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [18]),
        .Q(\main_inst/main_15_19_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [19]),
        .Q(\main_inst/main_15_19_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [20]),
        .Q(\main_inst/main_15_19_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [21]),
        .Q(\main_inst/main_15_19_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [22]),
        .Q(\main_inst/main_15_19_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [23]),
        .Q(\main_inst/main_15_19_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [24]),
        .Q(\main_inst/main_15_19_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [25]),
        .Q(\main_inst/main_15_19_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [26]),
        .Q(\main_inst/main_15_19_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [27]),
        .Q(\main_inst/main_15_19_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [28]),
        .Q(\main_inst/main_15_19_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [29]),
        .Q(\main_inst/main_15_19_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [30]),
        .Q(\main_inst/main_15_19_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [31]),
        .Q(\main_inst/main_15_19_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [32]),
        .Q(\main_inst/main_15_19_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [33]),
        .Q(\main_inst/main_15_19_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [34]),
        .Q(\main_inst/main_15_19_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [35]),
        .Q(\main_inst/main_15_19_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [36]),
        .Q(\main_inst/main_15_19_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [37]),
        .Q(\main_inst/main_15_19_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [38]),
        .Q(\main_inst/main_15_19_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [39]),
        .Q(\main_inst/main_15_19_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [40]),
        .Q(\main_inst/main_15_19_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [41]),
        .Q(\main_inst/main_15_19_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_15_19_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_15_17_reg ),
        .D(\main_inst/main_103_107 [10]),
        .Q(\main_inst/main_15_19_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [10]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [11]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [12]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [13]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [14]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [15]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [16]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [17]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [18]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [19]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [20]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [21]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [22]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [23]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [24]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [25]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [26]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [27]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [28]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [29]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [30]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [31]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [32]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [33]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [34]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [35]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [36]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [37]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [38]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [39]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [40]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_172_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_inst/main_103_107_reg [41]),
        .Q(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_169_expDiff1ii_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_169_expDiff1ii_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_169_expDiff1ii_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_169_expDiff1ii_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_169_expDiff1ii_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_169_172_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_169_expDiff1ii_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_ ),
        .Q(\main_inst/main_191_192_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[11] ),
        .Q(\main_inst/main_191_192_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[12] ),
        .Q(\main_inst/main_191_192_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[13] ),
        .Q(\main_inst/main_191_192_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[14] ),
        .Q(\main_inst/main_191_192_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[15] ),
        .Q(\main_inst/main_191_192_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[16] ),
        .Q(\main_inst/main_191_192_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[17] ),
        .Q(\main_inst/main_191_192_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[18] ),
        .Q(\main_inst/main_191_192_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[19] ),
        .Q(\main_inst/main_191_192_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[20] ),
        .Q(\main_inst/main_191_192_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[21] ),
        .Q(\main_inst/main_191_192_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[22] ),
        .Q(\main_inst/main_191_192_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[23] ),
        .Q(\main_inst/main_191_192_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[24] ),
        .Q(\main_inst/main_191_192_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[25] ),
        .Q(\main_inst/main_191_192_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[26] ),
        .Q(\main_inst/main_191_192_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[27] ),
        .Q(\main_inst/main_191_192_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[28] ),
        .Q(\main_inst/main_191_192_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[29] ),
        .Q(\main_inst/main_191_192_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[30] ),
        .Q(\main_inst/main_191_192_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[31] ),
        .Q(\main_inst/main_191_192_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[32] ),
        .Q(\main_inst/main_191_192_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[33] ),
        .Q(\main_inst/main_191_192_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[34] ),
        .Q(\main_inst/main_191_192_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[35] ),
        .Q(\main_inst/main_191_192_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[36] ),
        .Q(\main_inst/main_191_192_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[37] ),
        .Q(\main_inst/main_191_192_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[38] ),
        .Q(\main_inst/main_191_192_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[39] ),
        .Q(\main_inst/main_191_192_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[40] ),
        .Q(\main_inst/main_191_192_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_103_105_reg_reg_n_0_[41] ),
        .Q(\main_inst/main_191_192_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_192_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_192 ),
        .Q(\main_inst/main_191_192_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(main_191_193_reg),
        .Q(\main_inst/main_191_193_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [10]),
        .Q(\main_inst/main_191_193_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [11]),
        .Q(\main_inst/main_191_193_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [12]),
        .Q(\main_inst/main_191_193_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [13]),
        .Q(\main_inst/main_191_193_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [14]),
        .Q(\main_inst/main_191_193_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [15]),
        .Q(\main_inst/main_191_193_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [16]),
        .Q(\main_inst/main_191_193_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [17]),
        .Q(\main_inst/main_191_193_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [18]),
        .Q(\main_inst/main_191_193_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [19]),
        .Q(\main_inst/main_191_193_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [20]),
        .Q(\main_inst/main_191_193_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [21]),
        .Q(\main_inst/main_191_193_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [22]),
        .Q(\main_inst/main_191_193_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [23]),
        .Q(\main_inst/main_191_193_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [24]),
        .Q(\main_inst/main_191_193_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [25]),
        .Q(\main_inst/main_191_193_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [26]),
        .Q(\main_inst/main_191_193_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [27]),
        .Q(\main_inst/main_191_193_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [28]),
        .Q(\main_inst/main_191_193_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [29]),
        .Q(\main_inst/main_191_193_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [30]),
        .Q(\main_inst/main_191_193_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [31]),
        .Q(\main_inst/main_191_193_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [32]),
        .Q(\main_inst/main_191_193_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [33]),
        .Q(\main_inst/main_191_193_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [34]),
        .Q(\main_inst/main_191_193_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [35]),
        .Q(\main_inst/main_191_193_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [36]),
        .Q(\main_inst/main_191_193_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [37]),
        .Q(\main_inst/main_191_193_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [38]),
        .Q(\main_inst/main_191_193_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [39]),
        .Q(\main_inst/main_191_193_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [40]),
        .Q(\main_inst/main_191_193_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_inst/main_191_193 [41]),
        .Q(\main_inst/main_191_193_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_193_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(\main_191_193_reg[9]_i_1_n_0 ),
        .Q(\main_inst/main_191_193_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_191_aExp1ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_191_aExp1ii_reg ),
        .D(main_191_aExp1ii_reg),
        .Q(\main_inst/main_191_aExp1ii_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_0ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(main_195_0ii_reg),
        .Q(\main_inst/main_195_0ii_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \main_inst/main_195_196_reg[0]_i_1 
       (.I0(\main_inst/main_195_zExp0ii_reg ),
        .O(\main_inst/main_195_196 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [0]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [10]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [1]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [2]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [31]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_inst/main_195_196_reg_reg[31]_i_1 
       (.CI(\main_inst/main_195_196_reg_reg[8]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\main_inst/main_195_196_reg_reg[31]_i_1_n_4 ,\main_inst/main_195_196 [31],\main_inst/main_195_196 [10:9]}),
        .S({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [3]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [4]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_inst/main_195_196_reg_reg[4]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(\main_inst/main_195_196_reg_reg ),
        .CYINIT(\main_inst/main_195_zExp0ii_reg ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_195_196 [4:1]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [5]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [6]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [7]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [8]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_inst/main_195_196_reg_reg[8]_i_1 
       (.CI(\main_inst/main_195_196_reg_reg [3]),
        .CO({\main_inst/main_195_196_reg_reg[8]_i_1_n_0 ,\main_inst/main_195_196_reg_reg[8]_i_1_n_1 ,\main_inst/main_195_196_reg_reg[8]_i_1_n_2 ,\main_inst/main_195_196_reg_reg[8]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/main_195_196 [8:5]),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_196_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_196 [9]),
        .Q(\main_inst/main_195_196_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_197_reg_reg 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_197 ),
        .Q(\main_inst/main_195_197_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_199_reg_reg 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_199 ),
        .Q(\main_inst/main_195_iiiii ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [24]),
        .Q(\main_inst/main_195_200_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [25]),
        .Q(\main_inst/main_195_200_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [26]),
        .Q(\main_inst/main_195_200_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [27]),
        .Q(\main_inst/main_195_200_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [28]),
        .Q(\main_inst/main_195_200_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [29]),
        .Q(\main_inst/main_195_200_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [30]),
        .Q(\main_inst/main_195_200_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_200_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_200 [31]),
        .Q(\main_inst/main_195_200_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [24]),
        .Q(\main_inst/main_195_extracttiiii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [25]),
        .Q(\main_inst/main_195_extracttiiii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [26]),
        .Q(\main_inst/main_195_extracttiiii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [27]),
        .Q(\main_inst/main_195_extracttiiii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [28]),
        .Q(\main_inst/main_195_extracttiiii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [29]),
        .Q(\main_inst/main_195_extracttiiii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [30]),
        .Q(\main_inst/main_195_extracttiiii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_extracttiiii_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_195_196_reg ),
        .D(\main_inst/main_195_asinkiiii [31]),
        .Q(\main_inst/main_195_extracttiiii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_iiiii_reg_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(main_195_iiiii_reg),
        .Q(\main_inst/main_195_iiiii_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zExp0ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zExp0ii ),
        .Q(\main_inst/main_195_zExp0ii_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [0]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [10]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [11]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [12]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [13]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [14]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [15]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [16]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [17]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [18]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [19]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [1]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [20]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [21]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [22]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [23]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [24]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [25]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [26]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [27]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [28]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [29]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [2]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [30]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [31]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [32]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [33]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [34]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [35]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [36]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [37]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [38]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [39]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [3]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [40]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [41]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [42]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [43]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [44]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [45]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [46]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [47]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [48]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [49]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [4]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [50]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [51]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [52]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [53]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [54]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [55]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [56]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [57]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [58]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [59]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [5]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [60]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [61]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [62]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [63]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [6]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [7]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [8]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_195_zSig0ii_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_195_zSig0ii_reg ),
        .D(\main_inst/main_195_zSig0ii [9]),
        .Q(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_ ),
        .Q(\main_inst/main_1_scevgep_reg1 [3]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[10] ),
        .Q(\main_inst/main_1_scevgep_reg1 [13]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[11] ),
        .Q(\main_inst/main_1_scevgep_reg1 [14]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[12] ),
        .Q(\main_inst/main_1_scevgep_reg1 [15]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[13] ),
        .Q(\main_inst/main_1_scevgep_reg1 [16]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[14] ),
        .Q(\main_inst/main_1_scevgep_reg1 [17]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[15] ),
        .Q(\main_inst/main_1_scevgep_reg1 [18]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[16] ),
        .Q(\main_inst/main_1_scevgep_reg1 [19]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[17] ),
        .Q(\main_inst/main_1_scevgep_reg1 [20]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[18] ),
        .Q(\main_inst/main_1_scevgep_reg1 [21]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[19] ),
        .Q(\main_inst/main_1_scevgep_reg1 [22]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[1] ),
        .Q(\main_inst/main_1_scevgep_reg1 [4]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[20] ),
        .Q(\main_inst/main_1_scevgep_reg1 [23]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[21] ),
        .Q(\main_inst/main_1_scevgep_reg1 [24]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[22] ),
        .Q(\main_inst/main_1_scevgep_reg1 [25]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[23] ),
        .Q(\main_inst/main_1_scevgep_reg1 [26]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[24] ),
        .Q(\main_inst/main_1_scevgep_reg1 [27]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[25] ),
        .Q(\main_inst/main_1_scevgep_reg1 [28]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[26] ),
        .Q(\main_inst/main_1_scevgep_reg1 [29]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[27] ),
        .Q(\main_inst/main_1_scevgep_reg1 [30]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[28] ),
        .Q(\main_inst/main_1_scevgep_reg1 [31]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[29] ),
        .Q(\main_inst/main_1_2_reg_reg_n_0_ ),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[2] ),
        .Q(\main_inst/main_1_scevgep_reg1 [5]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[30] ),
        .Q(\main_inst/main_1_2_reg_reg_n_0_[30] ),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[31] ),
        .Q(\main_inst/main_1_2_reg_reg_n_0_[31] ),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[3] ),
        .Q(\main_inst/main_1_scevgep_reg1 [6]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[4] ),
        .Q(\main_inst/main_1_scevgep_reg1 [7]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[5] ),
        .Q(\main_inst/main_1_scevgep_reg1 [8]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[6] ),
        .Q(\main_inst/main_1_scevgep_reg1 [9]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[7] ),
        .Q(\main_inst/main_1_scevgep_reg1 [10]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[8] ),
        .Q(\main_inst/main_1_scevgep_reg1 [11]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_2_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_inst/main_float64_addexit_220_reg_reg_n_0_[9] ),
        .Q(\main_inst/main_1_scevgep_reg1 [12]),
        .R(main_1_2_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[0]),
        .Q(\main_inst/main_15_17 [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[10]),
        .Q(\main_inst/main_15_17 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[11]),
        .Q(\main_inst/main_15_17 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[12]),
        .Q(\main_inst/main_15_17 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[13]),
        .Q(\main_inst/main_15_17 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[14]),
        .Q(\main_inst/main_15_17 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[15]),
        .Q(\main_inst/main_15_17 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[16]),
        .Q(\main_inst/main_15_17 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[17]),
        .Q(\main_inst/main_15_17 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[18]),
        .Q(\main_inst/main_15_17 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[19]),
        .Q(\main_inst/main_15_17 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[1]),
        .Q(\main_inst/main_15_17 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[20]),
        .Q(\main_inst/main_15_17 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[21]),
        .Q(\main_inst/main_15_17 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[22]),
        .Q(\main_inst/main_15_17 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[23]),
        .Q(\main_inst/main_15_17 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[24]),
        .Q(\main_inst/main_15_17 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[25]),
        .Q(\main_inst/main_15_17 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[26]),
        .Q(\main_inst/main_15_17 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[27]),
        .Q(\main_inst/main_15_17 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[28]),
        .Q(\main_inst/main_15_17 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[29]),
        .Q(\main_inst/main_15_17 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[2]),
        .Q(\main_inst/main_15_17 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[30]),
        .Q(\main_inst/main_15_17 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[31]),
        .Q(\main_inst/main_15_17 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[3]),
        .Q(\main_inst/main_15_17 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[4]),
        .Q(\main_inst/main_15_17 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[5]),
        .Q(\main_inst/main_15_17 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[6]),
        .Q(\main_inst/main_15_17 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[7]),
        .Q(\main_inst/main_15_17 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[8]),
        .Q(\main_inst/main_15_17 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_3_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_a[9]),
        .Q(\main_inst/main_15_17 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[0]),
        .Q(\main_inst/main_103_107 [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[10]),
        .Q(\main_inst/main_103_107 [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[11]),
        .Q(\main_inst/main_103_107 [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[12]),
        .Q(\main_inst/main_103_107 [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[13]),
        .Q(\main_inst/main_103_107 [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[14]),
        .Q(\main_inst/main_103_107 [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[15]),
        .Q(\main_inst/main_103_107 [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[16]),
        .Q(\main_inst/main_103_107 [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[17]),
        .Q(\main_inst/main_103_107 [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[18]),
        .Q(\main_inst/main_103_107 [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[19]),
        .Q(\main_inst/main_103_107 [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[1]),
        .Q(\main_inst/main_103_107 [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[20]),
        .Q(\main_inst/main_103_107 [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[21]),
        .Q(\main_inst/main_103_107 [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[22]),
        .Q(\main_inst/main_103_107 [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[23]),
        .Q(\main_inst/main_103_107 [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[24]),
        .Q(\main_inst/main_103_107 [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[25]),
        .Q(\main_inst/main_103_107 [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[26]),
        .Q(\main_inst/main_103_107 [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[27]),
        .Q(\main_inst/main_103_107 [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[28]),
        .Q(\main_inst/main_103_107 [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[29]),
        .Q(\main_inst/main_103_107 [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[2]),
        .Q(\main_inst/main_103_107 [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[30]),
        .Q(\main_inst/main_103_107 [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[31]),
        .Q(\main_inst/main_103_107 [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[3]),
        .Q(\main_inst/main_103_107 [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[4]),
        .Q(\main_inst/main_103_107 [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[5]),
        .Q(\main_inst/main_103_107 [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[6]),
        .Q(\main_inst/main_103_107 [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[7]),
        .Q(\main_inst/main_103_107 [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[8]),
        .Q(\main_inst/main_103_107 [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_4_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_1_3_reg ),
        .D(memory_controller_out_b[9]),
        .Q(\main_inst/main_103_107 [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[0]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[8]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[8]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[12]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[12]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[12]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[12]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[16]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[16]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[16]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[16]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[0]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[20]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[20]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[20]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[20]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[24]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[24]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[24]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[24]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[28]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[28]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[0]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[28]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[28]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[0]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[4]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[4]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[4]_i_1_n_5 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[4]_i_1_n_4 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[8]_i_1_n_7 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_main_result02_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_1_2_reg ),
        .D(\main_1_main_result02_reg_reg[8]_i_1_n_6 ),
        .Q(\main_inst/main_1_main_result02_reg_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [23]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [24]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [25]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [26]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [27]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [28]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [29]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [30]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_1_scevgep_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_1_scevgep_reg ),
        .D(\main_inst/main_1_scevgep [31]),
        .Q(\main_inst/main_1_scevgep_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [10]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [11]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [12]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [13]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [14]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [15]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [16]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [17]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [18]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [19]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [20]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [21]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [22]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [23]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [24]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [25]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [26]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [27]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [28]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [29]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [30]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [31]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [32]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [33]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [34]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [35]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [36]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [37]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [38]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [39]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [40]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_30_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_inst/main_15_19_reg [9]),
        .Q(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_27_expDiff0i2i_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_27_expDiff0i2i_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[15]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[19]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[23]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[27]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[31]_i_2_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[3]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(\main_169_expDiff1ii_reg_reg[7]_i_1_VCC_1 ),
        .Q(\main_inst/main_27_expDiff0i2i_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_27_expDiff0i2i_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_27_expDiff0i2i_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_27_30_reg ),
        .D(main_169_expDiff1ii_reg_reg),
        .Q(\main_inst/main_27_expDiff0i2i_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [10]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [11]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [12]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [13]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [14]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [15]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [16]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [17]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [18]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [19]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [20]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [21]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [22]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [23]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [24]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [25]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [26]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [27]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [28]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [29]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [30]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [31]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [32]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [33]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [34]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [35]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [36]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [37]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [38]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [39]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [40]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_62_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(\main_inst/main_91_92 [9]),
        .Q(\main_inst/main_59_62_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_64_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(ONE_10),
        .Q(\main_inst/main_59_64_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_64_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(ONE_8),
        .Q(\main_inst/main_59_64_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_64_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(ONE_7),
        .Q(\main_inst/main_59_64_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_64_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(ONE_12),
        .Q(\main_inst/main_59_64_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_64_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(ONE_11),
        .Q(\main_inst/main_59_64_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_59_expDiff1i3i_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_59_62_reg ),
        .D(main_136_expDiff0ii_reg_reg),
        .Q(\main_inst/main_59_expDiff1i3i_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(main_float64_addexit_0i_reg),
        .Q(\main_inst/main_float64_addexit_0i_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[10]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[11]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[12]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[13]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[14]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[15]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[16]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[17]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[18]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[19]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[20]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[21]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[22]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[23]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[24]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[25]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[26]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[27]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[28]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[29]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[30]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[31]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[32]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[33]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[34]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[35]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[36]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[37]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[38]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[39]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[40]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[41]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[42]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[43]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[44]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[45]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[46]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[47]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[48]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[49]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[50]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[51]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[52]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[53]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[54]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[55]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[56]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[57]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[58]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[59]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[60]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[61]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[62]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[63]_inv 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[63]_inv_i_2_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_0i_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_0i_reg0 ),
        .D(\main_float64_addexit_0i_reg[9]_i_1_n_0 ),
        .Q(\main_inst/main_float64_addexit_0i_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [0]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [10]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [11]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [12]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [13]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [14]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [15]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [16]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [17]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [18]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [19]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [1]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [20]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [21]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [22]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [23]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [24]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [25]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [26]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [27]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [28]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [29]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [2]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [30]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [31]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [3]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [4]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [5]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [6]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [7]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [8]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_218_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_218_reg ),
        .D(\main_inst/main_float64_addexit_218 [9]),
        .Q(\main_inst/main_float64_addexit_218_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [0]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [10]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [11]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [12]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [13]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [14]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [15]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [16]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [17]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [18]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [19]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [1]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [20]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [21]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [22]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [23]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [24]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [25]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [26]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [27]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [28]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [29]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [2]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [30]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [31]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [3]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [4]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [5]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [6]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [7]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [8]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_220_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_220 [9]),
        .Q(\main_inst/main_float64_addexit_220_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_float64_addexit_exitcond1_reg_reg 
       (.C(clk),
        .CE(\main_inst/main_float64_addexit_220_reg ),
        .D(\main_inst/main_float64_addexit_exitcond1 ),
        .Q(\main_inst/main_float64_addexit_exitcond1_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ),
        .D(main_normalizeRoundAndPackFloat64exitii_209_reg),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ),
        .D(\main_inst/main_normalizeRoundAndPackFloat64exitii_209 ),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ),
        .D(\main_normalizeRoundAndPackFloat64exitii_209_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ),
        .D(\main_normalizeRoundAndPackFloat64exitii_209_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [0]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [10]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [11]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [12]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [13]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [14]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [15]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [16]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [17]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [18]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [19]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [1]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [20]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [21]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [22]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [23]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [24]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [25]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [26]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [27]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [28]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [29]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [2]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [30]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [31]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [32]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [33]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [34]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [35]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [36]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [37]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [38]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [39]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [3]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [40]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [41]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [42]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [43]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [44]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [45]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [46]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [47]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [48]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [49]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [4]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [50]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [51]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [52]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [53]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [54]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [55]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [56]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [57]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [58]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [59]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [5]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [60]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [61]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [62]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [63]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [6]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [7]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [8]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .D(\main_inst/roundAndPackFloat64_return_val_reg [9]),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[10] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [10]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[11] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [11]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[12] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [12]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[13] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [13]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[14] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [14]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[15] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [15]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[16] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [16]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[17] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [17]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[18] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [18]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[19] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [19]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[1] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [1]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[20] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [20]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[21] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [21]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[22] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [22]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[23] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [23]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[24] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [24]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[25] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [25]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[26] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [26]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[27] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [27]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[28] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [28]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[29] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [29]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[2] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [2]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[30] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [30]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[31] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [31]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[32] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [32]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[33] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [33]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[34] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [34]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[35] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [35]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[36] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [36]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[37] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [37]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[38] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [38]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[39] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [39]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[3] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [3]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[40] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [40]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[41] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [41]),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[4] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [4]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[5] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [5]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[6] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [6]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[7] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [7]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[8] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [8]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg_reg[9] 
       (.C(clk),
        .CE(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit3ii_z0i2ii_reg [9]),
        .R(ZERO_237));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_100_reg_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(main_shift64RightJammingexit9ii_100_reg),
        .Q(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[0]_i_1_n_0 ),
        .Q(\main_inst/A [0]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[10]_i_1_n_0 ),
        .Q(\main_inst/A [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[11]_i_1_n_0 ),
        .Q(\main_inst/A [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[12]_i_1_n_0 ),
        .Q(\main_inst/A [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[13]_i_1_n_0 ),
        .Q(\main_inst/A [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[14]_i_1_n_0 ),
        .Q(\main_inst/A [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[15]_i_1_n_0 ),
        .Q(\main_inst/A [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[16]_i_1_n_0 ),
        .Q(\main_inst/A [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[17]_i_1_n_0 ),
        .Q(\main_inst/A [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[18]_i_1_n_0 ),
        .Q(\main_inst/A [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[19]_i_1_n_0 ),
        .Q(\main_inst/A [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[1]_i_1_n_0 ),
        .Q(\main_inst/A [1]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[20]_i_1_n_0 ),
        .Q(\main_inst/A [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[21]_i_1_n_0 ),
        .Q(\main_inst/A [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[22]_i_1_n_0 ),
        .Q(\main_inst/A [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[23]_i_1_n_0 ),
        .Q(\main_inst/A [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[24]_i_1_n_0 ),
        .Q(\main_inst/A [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[25]_i_1_n_0 ),
        .Q(\main_inst/A [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[26]_i_1_n_0 ),
        .Q(\main_inst/A [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[27]_i_1_n_0 ),
        .Q(\main_inst/A [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[28]_i_1_n_0 ),
        .Q(\main_inst/A [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[29]_i_1_n_0 ),
        .Q(\main_inst/A [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[2]_i_1_n_0 ),
        .Q(\main_inst/A [2]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[30]_i_1_n_0 ),
        .Q(\main_inst/A [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[31]_i_1_n_0 ),
        .Q(\main_inst/A [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[32]_i_1_n_0 ),
        .Q(\main_inst/A [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[33]_i_1_n_0 ),
        .Q(\main_inst/A [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[34]_i_1_n_0 ),
        .Q(\main_inst/A [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[35]_i_1_n_0 ),
        .Q(\main_inst/A [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[36]_i_1_n_0 ),
        .Q(\main_inst/A [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[37]_i_1_n_0 ),
        .Q(\main_inst/A [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[38]_i_1_n_0 ),
        .Q(\main_inst/A [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[39]_i_1_n_0 ),
        .Q(\main_inst/A [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[3]_i_1_n_0 ),
        .Q(\main_inst/A [3]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[40]_i_1_n_0 ),
        .Q(\main_inst/A [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[4]_i_1_n_0 ),
        .Q(\main_inst/A [4]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[5]_i_1_n_0 ),
        .Q(\main_inst/A [5]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[6]_i_1_n_0 ),
        .Q(\main_inst/A [6]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[7]_i_1_n_0 ),
        .Q(\main_inst/A [7]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[8]_i_2_n_0 ),
        .Q(\main_inst/A [8]),
        .R(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_94_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_94_reg[9]_i_1_n_0 ),
        .Q(\main_inst/A [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[0]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[10]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[11]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[12]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[13]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[14]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[15]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[16]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[17]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[18]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[19]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[20]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[21]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[22]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[23]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[24]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[25]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[26]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[27]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[28]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[29]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[30]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[31]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[32]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[33]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[34]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[35]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[36]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[37]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[38]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[39]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_inst/main_shift64RightJammingexit9ii_95 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_95_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .D(\main_shift64RightJammingexit9ii_95_reg[9]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_95_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[63]_i_1_VCC_1 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_5 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_4 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_7 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexit9ii_ii_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/main_shift64RightJammingexit9ii_99_reg ),
        .D(\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_6 ),
        .Q(\main_inst/main_shift64RightJammingexit9ii_ii_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[0] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[0]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[10] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [10]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[11] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [11]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[12] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [12]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[13] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [13]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[14] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [14]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[15] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [15]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[16] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [16]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[17] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [17]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[18] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [18]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[19] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [19]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[1] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[1]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [1]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[20] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [20]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[21] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [21]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[22] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [22]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[23] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [23]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[24] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [24]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[25] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [25]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[26] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [26]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[27] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [27]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[28] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [28]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[29] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [29]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[2] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[2]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [2]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[30] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [30]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[31] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [31]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[32] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [32]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[33] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [33]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[34] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [34]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[35] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [35]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[36] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [36]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[37] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [37]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[38] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [38]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[39] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [39]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[3] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[3]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [3]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[40] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [40]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[41] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_inst/main_shift64RightJammingexitii_z0iii [41]),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[4] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[4]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [4]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[5] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[5]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [5]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[6] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[6]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [6]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[7] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[7]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [7]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[8] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[8]_i_1_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [8]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/main_shift64RightJammingexitii_z0iii_reg_reg[9] 
       (.C(clk),
        .CE(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ),
        .D(\main_shift64RightJammingexitii_z0iii_reg[9]_i_2_n_0 ),
        .Q(\main_inst/main_shift64RightJammingexitii_z0iii_reg [9]),
        .R(ZERO_245));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[0] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_ ),
        .Q(return_val[0]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[10] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[10] ),
        .Q(return_val[10]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[11] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[11] ),
        .Q(return_val[11]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[12] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[12] ),
        .Q(return_val[12]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[13] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[13] ),
        .Q(return_val[13]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[14] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[14] ),
        .Q(return_val[14]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[15] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[15] ),
        .Q(return_val[15]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[16] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[16] ),
        .Q(return_val[16]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[17] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[17] ),
        .Q(return_val[17]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[18] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[18] ),
        .Q(return_val[18]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[19] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[19] ),
        .Q(return_val[19]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[1] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[1] ),
        .Q(return_val[1]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[20] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[20] ),
        .Q(return_val[20]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[21] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[21] ),
        .Q(return_val[21]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[22] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[22] ),
        .Q(return_val[22]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[23] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[23] ),
        .Q(return_val[23]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[24] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[24] ),
        .Q(return_val[24]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[25] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[25] ),
        .Q(return_val[25]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[26] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[26] ),
        .Q(return_val[26]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[27] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[27] ),
        .Q(return_val[27]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[28] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[28] ),
        .Q(return_val[28]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[29] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[29] ),
        .Q(return_val[29]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[2] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[2] ),
        .Q(return_val[2]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[30] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[30] ),
        .Q(return_val[30]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[31] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[31] ),
        .Q(return_val[31]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[3] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[3] ),
        .Q(return_val[3]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[4] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[4] ),
        .Q(return_val[4]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[5] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[5] ),
        .Q(return_val[5]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[6] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[6] ),
        .Q(return_val[6]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[7] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[7] ),
        .Q(return_val[7]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[8] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[8] ),
        .Q(return_val[8]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/return_val_reg[9] 
       (.C(clk),
        .CE(\return_val[31]_i_2_n_0 ),
        .D(\main_inst/main_float64_addexit_218_reg_reg_n_0_[9] ),
        .Q(return_val[9]),
        .R(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/FSM_sequential_cur_state_reg[0] 
       (.C(clk),
        .CE(\FSM_sequential_cur_state[4]_i_1_n_0 ),
        .D(FSM_sequential_cur_state),
        .Q(\main_inst/roundAndPackFloat64/cur_state [0]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/FSM_sequential_cur_state_reg[1] 
       (.C(clk),
        .CE(\FSM_sequential_cur_state[4]_i_1_n_0 ),
        .D(FSM_sequential_cur_state_reg),
        .Q(\main_inst/roundAndPackFloat64/cur_state [1]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/FSM_sequential_cur_state_reg[2] 
       (.C(clk),
        .CE(\FSM_sequential_cur_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_cur_state_reg[2]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/cur_state [2]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/FSM_sequential_cur_state_reg[3] 
       (.C(clk),
        .CE(\FSM_sequential_cur_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_cur_state[3]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/cur_state [3]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* KEEP = "yes" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/FSM_sequential_cur_state_reg[4] 
       (.C(clk),
        .CE(\FSM_sequential_cur_state[4]_i_1_n_0 ),
        .D(\FSM_sequential_cur_state[4]_i_2_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/cur_state [4]),
        .R(reset));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/finish_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\main_inst/finish_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64_finish ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[0] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [0]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_ ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[10] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [10]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[10] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[11] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [11]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[11] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[12] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [12]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[12] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[13] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [13]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[13] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[14] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [14]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[14] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[15] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [15]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[15] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[16] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [16]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[16] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[17] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [17]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[17] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[18] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [18]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[18] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[19] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [19]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[19] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[1] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [1]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[1] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[20] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [20]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[20] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[21] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [21]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[21] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[22] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [22]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[22] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[23] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [23]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[23] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[24] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [24]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[24] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[25] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [25]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[25] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[26] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [26]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[26] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[27] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [27]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[27] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[28] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [28]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[28] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[29] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [29]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[29] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[2] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [2]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[2] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[30] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [30]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[30] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[31] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [31]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[31] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[32] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [32]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[32] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[33] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [33]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[33] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[34] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [34]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[34] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[35] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [35]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[35] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[36] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [36]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[36] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[37] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [37]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[37] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[38] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [38]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[38] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[39] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [39]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[39] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[3] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [3]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[3] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[40] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [40]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[40] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[41] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [41]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[41] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[42] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [42]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[42] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[43] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [43]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[43] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[44] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [44]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[44] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[45] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [45]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[45] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[46] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [46]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[46] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[47] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [47]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[47] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[48] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [48]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[48] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[49] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [49]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[49] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[4] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [4]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[4] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[50] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [50]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[50] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[51] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [51]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[51] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[52] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [52]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[52] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[53] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [53]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[53] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[54] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [54]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[54] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[55] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [55]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[55] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[56] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [56]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[56] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[57] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [57]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[57] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[58] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [58]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[58] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[59] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [59]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[59] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[5] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [5]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[5] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[60] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [60]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[60] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[61] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [61]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[61] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[62] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [62]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[62] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[63] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [63]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[63] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[6] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [6]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[6] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[7] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [7]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[7] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[8] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [8]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[8] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/return_val_reg[9] 
       (.C(clk),
        .CE(\return_val[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [9]),
        .Q(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[9] ),
        .R(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_11_16_reg_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(roundAndPackFloat64_11_16_reg),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_11_16_reg ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[0] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [0]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [0]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[10] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [10]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [10]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[11] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [11]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[12] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [12]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [12]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[13] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [13]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [13]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[14] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [14]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [14]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[15] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [15]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [15]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[16] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [16]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [16]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[17] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [17]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [17]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[18] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [18]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [18]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[19] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [19]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [19]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[1] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [1]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [1]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[20] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [20]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [20]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[21] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [21]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [21]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[22] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [22]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [22]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[23] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [23]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [23]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[24] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [24]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [24]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[25] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [25]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [25]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[26] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [26]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [26]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[27] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [27]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [27]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[28] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [28]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [28]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[29] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [29]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [29]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[2] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [2]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [2]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[30] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [30]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [30]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[31] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [31]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [31]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[32] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [32]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [32]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[33] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [33]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [33]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[34] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [34]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [34]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[35] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [35]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [35]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[36] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [36]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [36]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[37] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [37]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [37]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[38] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [38]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [38]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[39] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [39]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [39]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[3] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [3]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [3]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[40] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [40]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [40]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[41] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [41]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [41]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[42] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [42]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [42]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[43] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [43]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [43]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[44] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [44]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [44]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[45] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [45]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [45]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[46] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [46]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [46]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[47] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [47]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [47]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[48] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [48]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [48]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[49] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [49]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [49]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[4] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [4]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [4]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[50] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [50]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [50]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[51] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [51]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [51]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[52] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(roundAndPackFloat64_57_0_reg),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[53] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_6 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[54] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_5 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[55] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_4 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[56] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_7 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[57] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_6 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[58] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_5 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[59] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_4 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[5] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [5]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [5]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[60] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_7 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[61] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_6 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[62] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_5 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[63] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_4 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[6] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [6]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [6]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[7] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [7]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [7]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[8] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [8]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg_reg[9] 
       (.C(clk),
        .CE(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_57_0_reg [9]),
        .R(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [0]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [1]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [2]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [3]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [4]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [5]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [6]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [7]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[10] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [10]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[11] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [11]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[12] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [12]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[13] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [13]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[14] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [14]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[15] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [15]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[16] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [16]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[17] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [17]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[18] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [18]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[19] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [19]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[1] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [1]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[20] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [20]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[21] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [21]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[22] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [22]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[23] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [23]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[24] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [24]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[25] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [25]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[26] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [26]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[27] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [27]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[28] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [28]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[29] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [29]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[2] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [2]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[30] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [30]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[31] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [31]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[32] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [32]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[33] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [33]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[34] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [34]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[35] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [35]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[36] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [36]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[37] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [37]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[38] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [38]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[39] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [39]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[3] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [3]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[40] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [40]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[41] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [41]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[42] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [42]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[43] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [43]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[44] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [44]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[45] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [45]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[46] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [46]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[47] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [47]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[48] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [48]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[49] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [49]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[4] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [4]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[50] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [50]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[51] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [51]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[52] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [52]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[53] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [53]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[54] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [54]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[55] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [55]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[56] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [56]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[57] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [57]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[58] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [58]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[59] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [59]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[5] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [5]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[60] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [60]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[61] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [61]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[62] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_3_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [62]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[63] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[6] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [6]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[7] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [7]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[8] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [8]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[9] 
       (.C(clk),
        .CE(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .D(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [9]),
        .R(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [0]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [52]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [10]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [62]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [63]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [1]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [53]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [2]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [54]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [3]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [55]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [4]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [56]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [5]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [57]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [6]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [58]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [7]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [59]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [60]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_028_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [61]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [20]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [21]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [22]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [23]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [24]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [25]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [26]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [27]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [28]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [29]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [30]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [31]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [32]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [33]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [34]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [35]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [36]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [37]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [38]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [39]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [12]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [40]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [41]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [42]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [43]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [44]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [45]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [46]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [47]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [48]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [49]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [13]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [50]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [51]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [52]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [53]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [54]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [55]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [56]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [57]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [58]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [59]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [14]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [60]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [61]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [62]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [63]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [15]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64_arg_zSign_reg_n_0_ ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [16]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [17]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [18]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [19]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [52]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [53]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [54]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [55]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [56]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [57]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [58]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [59]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [60]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [61]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [62]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op [63]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_ ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [0]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[1] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [1]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[2] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [2]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[3] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [3]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[4] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [4]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[5] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [5]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[6] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [6]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[7] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [7]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[8] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [8]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[9] ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [9]),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [10]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [12]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [13]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [14]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [15]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [16]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [17]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [18]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [19]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [20]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [21]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [22]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [23]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [24]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [25]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [26]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [27]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [28]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [29]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [30]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [31]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [32]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [33]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [34]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [35]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [36]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [37]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [38]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [39]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [40]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [41]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [42]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [43]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [44]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [45]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [46]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [47]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [48]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [49]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [50]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [51]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [52]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [53]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [54]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [55]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [56]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [57]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [58]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [59]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [60]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [61]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [62]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [63]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[8] ),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[9] ),
        .R(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(roundAndPackFloat64_thread_02_reg),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [0]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[10]_i_2_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [10]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02 [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02 [1]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[2]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [2]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[3]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [3]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[4]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [4]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[5]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [5]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[6]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [6]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[7]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [7]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[8]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [8]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\roundAndPackFloat64_thread_02_reg[9]_i_1_n_0 ),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02_reg [9]),
        .R(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [0]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [1]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [2]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [3]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [4]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [5]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [6]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [7]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [10]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [11]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[12] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [12]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[13] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [13]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[14] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [14]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[15] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [15]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[16] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [16]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[17] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [17]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[18] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [18]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[19] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [19]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[20] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [20]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[21] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [21]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[22] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [22]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[23] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [23]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[24] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [24]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[25] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [25]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[26] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [26]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[27] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [27]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[28] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [28]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[29] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [29]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[30] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [30]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[31] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [31]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[32] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [32]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[33] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [33]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[34] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [34]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[35] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [35]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[36] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [36]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[37] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [37]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[38] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [38]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[39] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [39]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[40] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [40]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[41] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [41]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[42] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [42]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[43] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [43]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[44] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [44]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[45] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [45]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[46] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [46]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[47] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [47]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[48] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [48]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[49] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [49]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[50] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [50]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[51] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [51]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[52] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [52]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[53] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [53]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[54] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [54]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[55] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [55]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[56] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [56]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[57] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [57]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[58] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [58]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[59] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [59]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[60] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [60]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[61] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [61]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[62] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [62]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[63] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [63]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [8]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ),
        .D(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [9]),
        .Q(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \main_inst/roundAndPackFloat64_57_0_reg[51]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_57_0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [0]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [10]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [11]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[12] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [12]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[13] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [13]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[14] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [14]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[15] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [15]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[16] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [16]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[17] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [17]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[18] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [18]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[19] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [19]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [1]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[20] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [20]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[21] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [21]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[22] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [22]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[23] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [23]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[24] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [24]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[25] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [25]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[26] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [26]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[27] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [27]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[28] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [28]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[29] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [29]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [2]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[30] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [30]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[31] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [31]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [3]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [4]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [5]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [6]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [7]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [8]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zExp_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zExp [9]),
        .Q(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [0]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[10] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [10]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[11] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [11]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[12] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [12]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[13] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [13]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[14] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [14]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[15] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [15]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[16] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [16]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[17] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [17]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[18] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [18]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[19] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [19]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[1] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [1]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[20] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [20]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[21] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [21]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[22] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [22]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[23] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [23]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[24] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [24]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[25] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [25]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[26] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [26]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[27] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [27]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[28] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [28]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[29] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [29]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[2] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [2]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[30] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [30]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[31] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [31]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[32] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [32]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[33] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [33]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[34] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [34]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[35] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [35]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[36] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [36]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[37] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [37]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[38] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [38]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[39] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [39]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[3] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [3]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[40] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [40]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[41] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [41]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[42] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [42]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[43] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [43]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[44] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [44]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[45] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [45]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[46] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [46]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[47] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [47]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[48] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [48]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[49] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [49]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[4] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [4]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[50] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [50]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[51] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [51]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[52] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [52]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[53] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [53]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[54] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [54]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[55] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [55]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[56] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [56]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[57] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [57]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[58] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [58]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[59] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [59]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[5] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [5]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[60] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [60]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[61] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [61]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[62] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [62]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[63] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [63]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[6] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [6]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[7] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [7]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[8] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [8]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSig_reg[9] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(\main_inst/roundAndPackFloat64_arg_zSig [9]),
        .Q(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_arg_zSign_reg[0] 
       (.C(clk),
        .CE(\main_inst/roundAndPackFloat64_arg_zSign ),
        .D(roundAndPackFloat64_arg_zSign),
        .Q(\main_inst/roundAndPackFloat64_arg_zSign_reg_n_0_ ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_finish_reg_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(roundAndPackFloat64_finish_reg_i_1_n_0),
        .Q(\main_inst/roundAndPackFloat64_finish_reg_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[0] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_ ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [0]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[10] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[10] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [10]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[11] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[11] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [11]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[12] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[12] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [12]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[13] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[13] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [13]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[14] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[14] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [14]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[15] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[15] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [15]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[16] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[16] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [16]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[17] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[17] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [17]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[18] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[18] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [18]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[19] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[19] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [19]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[1] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[1] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [1]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[20] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[20] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [20]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[21] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[21] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [21]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[22] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[22] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [22]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[23] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[23] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [23]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[24] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[24] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [24]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[25] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[25] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [25]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[26] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[26] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [26]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[27] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[27] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [27]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[28] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[28] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [28]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[29] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[29] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [29]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[2] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[2] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [2]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[30] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[30] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [30]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[31] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[31] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [31]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[32] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[32] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [32]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[33] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[33] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [33]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[34] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[34] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [34]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[35] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[35] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [35]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[36] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[36] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [36]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[37] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[37] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [37]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[38] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[38] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [38]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[39] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[39] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [39]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[3] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[3] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [3]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[40] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[40] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [40]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[41] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[41] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [41]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[42] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[42] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [42]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[43] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[43] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [43]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[44] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[44] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [44]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[45] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[45] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [45]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[46] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[46] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [46]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[47] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[47] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [47]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[48] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[48] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [48]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[49] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[49] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [49]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[4] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[4] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [4]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[50] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[50] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [50]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[51] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[51] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [51]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[52] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[52] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [52]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[53] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[53] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [53]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[54] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[54] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [54]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[55] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[55] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [55]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[56] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[56] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [56]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[57] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[57] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [57]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[58] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[58] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [58]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[59] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[59] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [59]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[5] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[5] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [5]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[60] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[60] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [60]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[61] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[61] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [61]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[62] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[62] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [62]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[63] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[63] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [63]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[6] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[6] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [6]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[7] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[7] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [7]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[8] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[8] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [8]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_return_val_reg_reg[9] 
       (.C(clk),
        .CE(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ),
        .D(\main_inst/roundAndPackFloat64/return_val_reg_n_0_[9] ),
        .Q(\main_inst/roundAndPackFloat64_return_val_reg [9]),
        .R(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \main_inst/roundAndPackFloat64_start_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(roundAndPackFloat64_start_i_1_n_0),
        .Q(\main_inst/roundAndPackFloat64_start_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \main_normalizeRoundAndPackFloat64exitii_209_reg[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ),
        .O(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_normalizeRoundAndPackFloat64exitii_209_reg[31]_i_2 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .I2(\main_inst/main_195_197_reg ),
        .O(main_normalizeRoundAndPackFloat64exitii_209_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \main_normalizeRoundAndPackFloat64exitii_209_reg[3]_i_1 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .O(\main_inst/main_normalizeRoundAndPackFloat64exitii_209 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair362" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \main_normalizeRoundAndPackFloat64exitii_209_reg[4]_i_1 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ),
        .O(\main_normalizeRoundAndPackFloat64exitii_209_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    \main_normalizeRoundAndPackFloat64exitii_209_reg[5]_i_1 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ),
        .I1(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .I2(\main_inst/main_195_197_reg ),
        .O(\main_normalizeRoundAndPackFloat64exitii_209_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \main_normalizeRoundAndPackFloat64exitii_214_reg[63]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\return_val[31]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00FF0040)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[3]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_1_2_reg[31]_i_4_n_0 ),
        .I3(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_3_n_0 ),
        .I4(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_ ),
        .O(main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAFCFFAAAA0C00)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_1 
       (.I0(\main_inst/main_195_iiiii ),
        .I1(\main_inst/main_195_iiiii_reg ),
        .I2(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ),
        .I3(\main_1_2_reg[31]_i_4_n_0 ),
        .I4(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_3_n_0 ),
        .I5(\main_inst/main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg_reg_n_0_[4] ),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000BFFF00000000)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_3 
       (.I0(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_4_n_0 ),
        .I1(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_5_n_0 ),
        .I2(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_6_n_0 ),
        .I3(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_7_n_0 ),
        .I4(\main_195_zSig0ii_reg[63]_i_3_n_0 ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFACFCA)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_4 
       (.I0(\main_inst/main_195_extracttiiii_reg [28]),
        .I1(\main_inst/main_195_200_reg [28]),
        .I2(\main_inst/main_195_iiiii ),
        .I3(\main_inst/main_195_extracttiiii_reg [29]),
        .I4(\main_inst/main_195_200_reg [29]),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053035)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_5 
       (.I0(\main_inst/main_195_extracttiiii_reg [31]),
        .I1(\main_inst/main_195_200_reg [31]),
        .I2(\main_inst/main_195_iiiii ),
        .I3(\main_inst/main_195_extracttiiii_reg [30]),
        .I4(\main_inst/main_195_200_reg [30]),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053035)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_6 
       (.I0(\main_inst/main_195_extracttiiii_reg [26]),
        .I1(\main_inst/main_195_200_reg [26]),
        .I2(\main_inst/main_195_iiiii ),
        .I3(\main_inst/main_195_extracttiiii_reg [27]),
        .I4(\main_inst/main_195_200_reg [27]),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00053035)) 
    \main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_7 
       (.I0(\main_inst/main_195_extracttiiii_reg [24]),
        .I1(\main_inst/main_195_200_reg [24]),
        .I2(\main_inst/main_195_iiiii ),
        .I3(\main_inst/main_195_extracttiiii_reg [25]),
        .I4(\main_inst/main_195_200_reg [25]),
        .O(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_10 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_7_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_100 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .O(main_shift64RightJammingexit3ii_z0i2ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_101 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_102 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_103 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_104 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[14] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_105 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[13] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[11] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h0D)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_106 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_136_expDiff0ii_reg ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_ ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_141 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_142 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[15] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_143 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[12] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_144 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_ ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[11] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEAEFFFFFEAE0000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_2 
       (.I0(\main_inst/main_145_152 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_4_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_2_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I5(\main_inst/main_154_156 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_27 
       (.I0(\main_inst/main_136_expDiff0ii_reg ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_28 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_29 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_30 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_4 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_3_n_0 ),
        .I3(\main_inst/main_136_141_reg [2]),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_58 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_59 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_60 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_62 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_63 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_64 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_65 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_136_expDiff0ii_reg ),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_99 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3_n_0 ),
        .I3(\main_inst/main_136_141_reg [1]),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[14] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_2_n_0 ),
        .I5(\main_inst/main_136_expDiff0ii_reg ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_3_n_0 ),
        .I3(\main_inst/main_136_141_reg [1]),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_7_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .I5(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[30] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ),
        .I2(\main_inst/main_136_141_reg [1]),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[27] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[28] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_3_n_0 ),
        .I4(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[29] ),
        .I4(\main_inst/main_136_141_reg [4]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_inst/main_136_expDiff0ii_reg ),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_6_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_3 
       (.I0(\main_inst/main_136_141_reg [4]),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_141_reg [3]),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[26]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_3 
       (.I0(\main_inst/main_136_141_reg [4]),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_141_reg [3]),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[27]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_3 
       (.I0(\main_inst/main_136_141_reg [4]),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_141_reg [3]),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[28]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_3 
       (.I0(\main_inst/main_136_141_reg [4]),
        .I1(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_141_reg [3]),
        .I4(\main_inst/main_136_141_reg [2]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[29]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_inst/main_136_141_reg [4]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_141_reg [3]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_inst/main_136_141_reg [4]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_141_reg [3]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_inst/main_136_141_reg [4]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_141_reg [3]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_3 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_inst/main_136_141_reg [4]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_141_reg [3]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_3 
       (.I0(\main_inst/main_136_141_reg [3]),
        .I1(\main_inst/main_136_141_reg [5]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [2]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_4 
       (.I0(\main_inst/main_136_141_reg [3]),
        .I1(\main_inst/main_136_141_reg [5]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [2]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_3 
       (.I0(\main_inst/main_136_141_reg [3]),
        .I1(\main_inst/main_136_141_reg [5]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [2]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_4 
       (.I0(\main_inst/main_136_141_reg [3]),
        .I1(\main_inst/main_136_141_reg [5]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [2]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_2_n_0 ),
        .I5(\main_inst/main_136_expDiff0ii_reg ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_2_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_5_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_2 
       (.I0(\main_inst/main_136_141_reg [2]),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hAB)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_inst/main_136_expDiff0ii_reg ),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_5_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit3ii_z0i2ii [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_158_160_reg[62]_i_4_n_0 ),
        .I5(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFBFFFFFFFFFF)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_5 
       (.I0(\main_inst/main_136_141_reg [2]),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_inst/main_136_expDiff0ii_reg ),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_5_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_2_n_0 ),
        .I5(\main_inst/main_136_expDiff0ii_reg ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_inst/main_136_expDiff0ii_reg ),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_2_n_0 ),
        .I5(\main_inst/main_136_expDiff0ii_reg ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_4_n_0 ),
        .I1(\main_inst/main_136_141_reg [3]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_136_141_reg [4]),
        .I4(\main_inst/main_136_141_reg [5]),
        .I5(\main_inst/main_136_139_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_1 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2_n_0 ),
        .I1(\main_inst/main_136_141_reg [1]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I4(\main_inst/main_136_expDiff0ii_reg ),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[14]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[12]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_4 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_5 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_7_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_6 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_ ),
        .I3(\main_inst/main_136_141_reg [5]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_7 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[40] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_2 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[41]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_4_n_0 ),
        .I2(\main_inst/main_136_expDiff0ii_reg ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[10]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_4 
       (.I0(\main_shift64RightJammingexit3ii_z0i2ii_reg[15]_i_3_n_0 ),
        .I1(\main_inst/main_136_141_reg [2]),
        .I2(\main_shift64RightJammingexit3ii_z0i2ii_reg[11]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit3ii_z0i2ii_reg[13]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ),
        .I5(\main_inst/main_136_141_reg [1]),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_139_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_136_141_reg [5]),
        .I4(\main_inst/main_136_141_reg [3]),
        .I5(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_7_n_0 ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_7 
       (.I0(\main_inst/main_136_139_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_136_141_reg [4]),
        .I2(\main_inst/main_136_141_reg [5]),
        .I3(\main_inst/main_136_139_reg_reg_n_0_[41] ),
        .O(\main_shift64RightJammingexit3ii_z0i2ii_reg[9]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_11 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_0 ),
        .CO(main_shift64RightJammingexit3ii_z0i2ii_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_27_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_28_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_29_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_25_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_58_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_59_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_60_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_26_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_62_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_63_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_64_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_65_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_0 ,\main_inst/main_145_152 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,ONE_28,ONE_21,ONE_20}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5 
       (.CI(main_shift64RightJammingexit3ii_z0i2ii_reg_reg[3]),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_1 ,\main_inst/main_154_156 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_57_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_99_n_0 ,main_shift64RightJammingexit3ii_z0i2ii_reg,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_101_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_102_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6 
       (.CI(\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_12_n_0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({ONE_25,ONE_24,ONE_23,ONE_22}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_61_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_103_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_104_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_105_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_106_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_1 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_2 ,\main_shift64RightJammingexit3ii_z0i2ii_reg_reg[0]_i_98_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_141_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_142_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_143_n_0 ,\main_shift64RightJammingexit3ii_z0i2ii_reg[0]_i_144_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFF0001)) 
    \main_shift64RightJammingexit9ii_100_reg[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_shift64RightJammingexit9ii_100_reg[0]_i_2_n_0 ),
        .I4(\main_inst/main_shift64RightJammingexit9ii_100_reg_reg_n_0_ ),
        .O(main_shift64RightJammingexit9ii_100_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h7FFF)) 
    \main_shift64RightJammingexit9ii_100_reg[0]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_shift64RightJammingexit9ii_100_reg[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hCA)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_2 ),
        .I1(\main_inst/main_68_76 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_107 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .O(main_shift64RightJammingexit9ii_94_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_108 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[14] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_109 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[13] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[14] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[11] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0051)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_110 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_ ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[11] ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[9] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_12 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_16_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_14 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_15 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_16 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEAE)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_3 
       (.I0(\main_inst/main_68_75 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[0]_i_6_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[1]_i_2_n_0 ),
        .O(\main_inst/main_68_76 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_31 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_32 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_33 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_34 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0111)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_37 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_38 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_39 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_6 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[2]_i_3_n_0 ),
        .I3(\main_inst/main_59_64_reg [1]),
        .I4(\main_shift64RightJammingexit9ii_94_reg[4]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_94_reg[0]_i_12_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_66 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_67 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[15] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_68 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[12] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_69 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_ ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[9] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_71 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_72 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_73 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_94_reg[0]_i_74 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[0]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[10]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[10]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [10]),
        .O(\main_shift64RightJammingexit9ii_94_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[10]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[10]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[11]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[10]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[14]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[6]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[11]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[11]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [11]),
        .O(\main_shift64RightJammingexit9ii_94_reg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[11]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[11]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[11]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[12]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[12]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [12]),
        .O(\main_shift64RightJammingexit9ii_94_reg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[12]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[13]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[12]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_5_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[13]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[13]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [13]),
        .O(\main_shift64RightJammingexit9ii_94_reg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[13]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[13]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[13]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[14]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[14]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [14]),
        .O(\main_shift64RightJammingexit9ii_94_reg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[14]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[15]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[14]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[18]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[14]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[14]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[6]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[15]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[15]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [15]),
        .O(\main_shift64RightJammingexit9ii_94_reg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[15]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[15]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[15]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [16]),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[16]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[17]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[18]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_4 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[20]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[16]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_5 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[16]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[16]_i_6 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[16]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[17]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[17]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [17]),
        .O(\main_shift64RightJammingexit9ii_94_reg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[17]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[17]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[18]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[17]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[17]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[18]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[18]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [18]),
        .O(\main_shift64RightJammingexit9ii_94_reg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[18]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[18]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[19]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[18]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[20]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[18]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[18]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[19]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[19]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [19]),
        .O(\main_shift64RightJammingexit9ii_94_reg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[19]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[19]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[20]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[19]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[19]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[1]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[2]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[1]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexit9ii_94_reg[1]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[3]_i_3_n_0 ),
        .I3(\main_inst/main_59_64_reg [1]),
        .I4(\main_shift64RightJammingexit9ii_94_reg[5]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_94_reg[1]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[1]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_14_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[20]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[20]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [20]),
        .O(\main_shift64RightJammingexit9ii_94_reg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[20]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[20]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[21]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[20]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[20]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[20]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[21]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[21]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [21]),
        .O(\main_shift64RightJammingexit9ii_94_reg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[21]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[21]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[22]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[21]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[21]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[22]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[22]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [22]),
        .O(\main_shift64RightJammingexit9ii_94_reg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[22]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[22]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[23]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[22]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[22]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[22]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[23]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[23]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [23]),
        .O(\main_shift64RightJammingexit9ii_94_reg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[23]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[23]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[24]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[23]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[29]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[23]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[24]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[24]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [24]),
        .O(\main_shift64RightJammingexit9ii_94_reg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[24]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[24]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[25]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[24]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[26]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_94_reg[24]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .I5(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[25]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[25]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [25]),
        .O(\main_shift64RightJammingexit9ii_94_reg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[25]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[25]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[26]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[25]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[31]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[29]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[25]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[26]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[26]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [26]),
        .O(\main_shift64RightJammingexit9ii_94_reg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[26]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[27]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[26]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_94_reg[26]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[28]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ),
        .I2(\main_inst/main_59_64_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_94_reg[26]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[26]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[26]_i_5 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[27]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[27]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [27]),
        .O(\main_shift64RightJammingexit9ii_94_reg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[27]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[27]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[28]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[27]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[31]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[27]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[28]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[28]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [28]),
        .O(\main_shift64RightJammingexit9ii_94_reg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[28]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[28]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit9ii_94_reg[28]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[28]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[30]_i_4_n_0 ),
        .I4(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[28]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[28]_i_5 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[29]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[29]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [29]),
        .O(\main_shift64RightJammingexit9ii_94_reg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[29]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[30]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_94_reg[29]_i_3 
       (.I0(\main_inst/main_59_64_reg [4]),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_64_reg [3]),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[29]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[29]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[2]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[3]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[2]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[2]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[4]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[2]_i_3_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[2]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[6]_i_5_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[30]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[30]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [30]),
        .O(\main_shift64RightJammingexit9ii_94_reg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[30]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[30]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[30]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[32]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[30]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_94_reg[30]_i_4 
       (.I0(\main_inst/main_59_64_reg [4]),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_64_reg [3]),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[26]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[31]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[31]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [31]),
        .O(\main_shift64RightJammingexit9ii_94_reg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[31]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[32]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_94_reg[31]_i_3 
       (.I0(\main_inst/main_59_64_reg [4]),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_64_reg [3]),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[31]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[31]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_59_64_reg [4]),
        .O(\main_shift64RightJammingexit9ii_94_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[32]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[32]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [32]),
        .O(\main_shift64RightJammingexit9ii_94_reg[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[32]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[32]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[32]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[34]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[32]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_94_reg[32]_i_4 
       (.I0(\main_inst/main_59_64_reg [4]),
        .I1(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_64_reg [3]),
        .I4(\main_inst/main_59_64_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[28]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[33]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[33]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [33]),
        .O(\main_shift64RightJammingexit9ii_94_reg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[33]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[34]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[33]_i_3 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_inst/main_59_64_reg [4]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_64_reg [3]),
        .O(\main_shift64RightJammingexit9ii_94_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[34]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[34]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [34]),
        .O(\main_shift64RightJammingexit9ii_94_reg[34]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[34]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[34]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[34]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[36]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[34]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[34]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_inst/main_59_64_reg [4]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_64_reg [3]),
        .O(\main_shift64RightJammingexit9ii_94_reg[34]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[35]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[35]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [35]),
        .O(\main_shift64RightJammingexit9ii_94_reg[35]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[35]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[36]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[35]_i_3 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_inst/main_59_64_reg [4]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_64_reg [3]),
        .O(\main_shift64RightJammingexit9ii_94_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[36]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[36]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [36]),
        .O(\main_shift64RightJammingexit9ii_94_reg[36]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[36]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[37]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[36]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[36]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[38]_i_5_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[36]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_94_reg[36]_i_4 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_inst/main_59_64_reg [4]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_64_reg [3]),
        .O(\main_shift64RightJammingexit9ii_94_reg[36]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[37]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[37]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [37]),
        .O(\main_shift64RightJammingexit9ii_94_reg[37]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFB800B800000000)) 
    \main_shift64RightJammingexit9ii_94_reg[37]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[37]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ),
        .I3(\main_inst/main_59_expDiff1i3i_reg ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[38]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_94_reg[37]_i_3 
       (.I0(\main_inst/main_59_64_reg [3]),
        .I1(\main_inst/main_59_64_reg [5]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [2]),
        .O(\main_shift64RightJammingexit9ii_94_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_94_reg[37]_i_4 
       (.I0(\main_inst/main_59_64_reg [3]),
        .I1(\main_inst/main_59_64_reg [5]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [2]),
        .O(\main_shift64RightJammingexit9ii_94_reg[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[38]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[38]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [38]),
        .O(\main_shift64RightJammingexit9ii_94_reg[38]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[38]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[38]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[39]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_94_reg[38]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[38]_i_4_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[38]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_94_reg[38]_i_4 
       (.I0(\main_inst/main_59_64_reg [3]),
        .I1(\main_inst/main_59_64_reg [5]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [2]),
        .O(\main_shift64RightJammingexit9ii_94_reg[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_94_reg[38]_i_5 
       (.I0(\main_inst/main_59_64_reg [3]),
        .I1(\main_inst/main_59_64_reg [5]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [2]),
        .O(\main_shift64RightJammingexit9ii_94_reg[38]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[39]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[39]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [39]),
        .O(\main_shift64RightJammingexit9ii_94_reg[39]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hE200)) 
    \main_shift64RightJammingexit9ii_94_reg[39]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[39]_i_3_n_0 ),
        .I1(\main_inst/main_59_expDiff1i3i_reg ),
        .I2(\main_shift64RightJammingexit9ii_94_reg[40]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit9ii_94_reg[39]_i_3 
       (.I0(\main_inst/main_59_64_reg [2]),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[3]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[4]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[3]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[3]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[5]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[3]_i_3_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[3]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_12_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[40]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[40]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [40]),
        .O(\main_shift64RightJammingexit9ii_94_reg[40]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \main_shift64RightJammingexit9ii_94_reg[40]_i_2 
       (.I0(\main_inst/main_59_expDiff1i3i_reg ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[40]_i_3_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit9ii_94_reg[40]_i_3 
       (.I0(\main_inst/main_59_64_reg [2]),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[40]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[4]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[5]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[4]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[4]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[6]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[4]_i_3_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[4]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_15_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[5]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[6]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[5]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[5]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[5]_i_3_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[5]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_13_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[7]_i_2_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[6]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_9_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[6]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_3 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[6]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_4 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[6]_i_6_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_5 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_ ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[6]_i_6 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[14] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[6]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[7]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[8]_i_4_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[7]_i_2_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[7]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_94_reg[7]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_11_n_0 ),
        .I1(\main_inst/main_59_64_reg [3]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_59_64_reg [4]),
        .I4(\main_inst/main_59_64_reg [5]),
        .I5(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE0)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I2(\main_inst/main_shift64RightJammingexit9ii_94_reg ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_10 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_16_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_11 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_12 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_13 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_14 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[9] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_15 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_16 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_64_reg [5]),
        .I3(\main_inst/main_59_62_reg_reg_n_0_[40] ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8A80)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_94_reg[8]_i_3_n_0 ),
        .I2(\main_inst/main_59_expDiff1i3i_reg ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ),
        .I5(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_4 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[8]_i_9_n_0 ),
        .I1(\main_inst/main_59_64_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[8]_i_10_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[10]_i_3_n_0 ),
        .I4(\main_inst/main_59_64_reg [1]),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_5 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_11_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_6 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_12_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_7 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_13_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_8 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_14_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_94_reg[8]_i_9 
       (.I0(\main_inst/main_59_62_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_59_64_reg [4]),
        .I2(\main_inst/main_59_62_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_59_64_reg [5]),
        .I4(\main_inst/main_59_64_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_94_reg[8]_i_15_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE02)) 
    \main_shift64RightJammingexit9ii_94_reg[9]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[9]_i_2_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I3(\main_inst/main_91_92 [9]),
        .O(\main_shift64RightJammingexit9ii_94_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8FF0000000000)) 
    \main_shift64RightJammingexit9ii_94_reg[9]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_94_reg[12]_i_3_n_0 ),
        .I1(\main_inst/main_59_64_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_94_reg[10]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_94_reg[8]_i_3_n_0 ),
        .I4(\main_inst/main_59_expDiff1i3i_reg ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_shift64RightJammingexit9ii_94_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_13 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_0 ),
        .CO(main_shift64RightJammingexit9ii_94_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_94_reg[0]_i_31_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_32_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_33_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_34_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({ONE_13,\main_shift64RightJammingexit9ii_94_reg[0]_i_37_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_38_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_39_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_30_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_94_reg[0]_i_66_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_67_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_68_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_69_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_35_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_94_reg[0]_i_71_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_72_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_73_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_74_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_0 ,\main_inst/main_68_75 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,ONE_27,ONE_19,ONE_18}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7 
       (.CI(main_shift64RightJammingexit9ii_94_reg_reg[3]),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_14_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_15_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_70_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({main_shift64RightJammingexit9ii_94_reg,\main_shift64RightJammingexit9ii_94_reg[0]_i_108_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_109_n_0 ,\main_shift64RightJammingexit9ii_94_reg[0]_i_110_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8 
       (.CI(\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_17_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_0 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_1 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_2 ,\main_shift64RightJammingexit9ii_94_reg_reg[0]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({ONE_17,ONE_16,ONE_15,ONE_14}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_1 
       (.I0(\main_inst/main_45_47 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I3(\main_inst/main_35_44 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_10 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_24_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_23_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_25_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_26_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_100 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(main_shift64RightJammingexit9ii_95_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_101 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_102 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_103 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_156_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_104 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_157_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_105 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_106 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_106_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_107 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_158_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_108 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_159_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_109 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_11 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_27_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_26_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_28_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_29_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_110 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_111 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_160_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_111_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_112 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_161_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_113 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_114 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_115 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_162_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_130_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_163_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_164_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_116 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_165_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_164_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_166_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_167_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_117 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_168_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_167_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_169_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_170_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h005FFFFFFFFFF0F1)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_118 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_171_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_172_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_173_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_119 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_174_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_119_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_12 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_19_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_120 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_175_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_120_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_121 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_174_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_121_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_122 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_175_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_122_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_123 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_178_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_123_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_124 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_179_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_124_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_125 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_180_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_178_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_125_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_126 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_181_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_179_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_126_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_127 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_180_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_182_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_127_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_128 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_181_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_183_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_128_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_129 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_182_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_184_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_129_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_130 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_183_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_185_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_130_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_131 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_186_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_131_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_132 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_153_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_187_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_132_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_133 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_154_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_137_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_133_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_134 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_188_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_135 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_131_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_189_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_135_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_136 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_187_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_190_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_136_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_137 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_191_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_137_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_138 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_139 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_14 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_140 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_189_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_192_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_140_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_141 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_190_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_193_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_142 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_143 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_144 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_194_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_145 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_195_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_145_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_146 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_146_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_147 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_147_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_148 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_148_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_149 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_196_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_149_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_15 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_150 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_197_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_150_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_151 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_151_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_152 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_152_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_153 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_198_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_153_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_154 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_199_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_154_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_155 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_155_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_156 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_156_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_157 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_157_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_158 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_158_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_159 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_159_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_16 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_160 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_160_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_161 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_161_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_162 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_184_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_200_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_162_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_163 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_185_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_201_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_163_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_164 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_200_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_202_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_164_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_165 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_201_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_203_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_165_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_166 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_202_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_204_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_166_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBE82828282828282)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_167 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_203_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_205_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_167_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBE82828282828282)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_168 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_204_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_206_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_168_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBC80000000000202)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_169 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_205_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_207_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_169_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBC80000000000202)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_170 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_206_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_208_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_170_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_171 
       (.I0(main_shift64RightJammingexit9ii_95_reg),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_171_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_172 
       (.I0(main_shift64RightJammingexit9ii_95_reg),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_172_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_173 
       (.I0(main_shift64RightJammingexit9ii_95_reg),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_173_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_174 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_192_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_209_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_174_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_175 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_193_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_210_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_175_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_176 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_176_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_177 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_177_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_178 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_209_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_211_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_178_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_179 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_210_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_212_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_179_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_18 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_40_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_29_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_41_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_42_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_180 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_180_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_181 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_181_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_182 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_211_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_213_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_182_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_183 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_212_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_183_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_184 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_180_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_184_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_185 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_181_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_185_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_186 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_186_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_187 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_215_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_187_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_188 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_188_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_189 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_216_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_189_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_19 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_43_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_42_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_44_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_45_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_190 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_190_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_191 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_191_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_192 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_192_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_193 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_193_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_194 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_194_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_195 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_195_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_196 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_196_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_197 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_197_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_198 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_198_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_199 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_199_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_20 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_46_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_45_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_47_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_48_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_200 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_213_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_200_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_201 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_201_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_202 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_202_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_203 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_203_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_204 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_204_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_205 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_205_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_206 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_206_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_207 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_207_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_208 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_208_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_209 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I2(main_shift64RightJammingexit9ii_95_reg),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_209_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_21 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_49_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_48_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_50_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_51_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0008000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_210 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_210_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_211 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_211_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_212 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_212_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_213 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I1(main_shift64RightJammingexit9ii_95_reg),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_213_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_214 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_214_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_215 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_215_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_216 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_216_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFE2B80000E2)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_22 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_52_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_53_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_54_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFE2B80000E2)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_23 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_55_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_56_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_57_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_24 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_53_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_54_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_25 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_56_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_57_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_26 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_53_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_60_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_27 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_56_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_61_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_28 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_62_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_60_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_29 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_61_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFEAE)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_3 
       (.I0(\main_inst/main_35_43 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_6_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[1]_i_2_n_0 ),
        .O(\main_inst/main_35_44 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_31 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_32 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_33 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_34 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_36 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_73_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_51_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_74_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_75_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_37 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_76_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_75_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_77_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_78_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_38 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_79_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_78_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_80_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_81_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_39 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_82_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_81_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_83_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_84_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_40 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_62_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_85_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_41 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_86_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_42 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_85_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_87_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_43 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_86_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_44 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_89_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_87_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_45 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_91_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_46 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_89_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_92_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_47 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_91_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_48 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_92_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_49 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_95_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_50 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_96_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_51 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_95_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_52 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_101_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_53 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_102_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_54 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_103_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_104_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_55 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_105_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_56 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_106_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_57 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_107_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_108_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_58 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_109_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_59 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_110_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_6 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[2]_i_3_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[4]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_12_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_60 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_104_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_111_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_61 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_108_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_112_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_62 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_113_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_63 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_114_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_64 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_65 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_66 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_67 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_69 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_119_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_84_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_120_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_121_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_70 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_122_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_121_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_123_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_124_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_71 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_125_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_124_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_126_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_127_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_72 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_128_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_127_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_129_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_130_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_73 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_131_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_96_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_74 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_132_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_75 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_131_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_133_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_76 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_132_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_77 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_133_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_135_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_78 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_136_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_79 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_137_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_135_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_80 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_136_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_81 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_137_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_140_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_82 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_134_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_141_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_83 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_138_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_142_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_140_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_84 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_139_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_143_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_141_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_85 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_111_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_86 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_112_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_144_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_87 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_62_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_145_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_88 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_146_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_89 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_147_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_9 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_22_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[0]_i_23_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_90 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_148_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_91 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_144_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_149_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_92 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_145_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_150_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_93 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_151_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_94 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_152_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_95 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_149_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_153_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_96 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[0]_i_150_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[0]_i_154_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_97 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ),
        .I4(main_shift64RightJammingexit9ii_95_reg),
        .I5(\main_shift64RightJammingexit9ii_95_reg[0]_i_155_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFE0001)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_98 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000001)) 
    \main_shift64RightJammingexit9ii_95_reg[0]_i_99 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[0]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[10]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[11]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[10]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [10]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[10]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[11]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[12]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[11]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [11]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[11]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[12]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[13]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[12]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [12]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[12]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[13]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[14]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[13]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [13]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[13]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[14]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[15]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[14]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [14]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[14]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[15]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[16]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[15]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [15]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[15]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[16]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[17]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[16]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [16]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[16]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[16]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[16]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[16]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[16]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[17]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[18]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[17]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [17]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[17]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[17]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[18]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[19]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[18]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [18]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[18]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[18]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[19]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[20]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[19]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [19]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[19]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[19]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[1]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[2]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[1]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexit9ii_95_reg[1]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[3]_i_3_n_0 ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[5]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[1]_i_3_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[1]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_15_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[20]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[21]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[20]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [20]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[20]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[20]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[21]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[22]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[21]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [21]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[21]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[21]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[22]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[23]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[22]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [22]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[22]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[22]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[22]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[23]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[24]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[23]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [23]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[23]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[25]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[23]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[24]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[25]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[24]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [24]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[24]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[26]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexit9ii_95_reg[24]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[25]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[26]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[25]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [25]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[25]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[27]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[25]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[25]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[25]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[25]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[26]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[27]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[26]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [26]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexit9ii_95_reg[26]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[28]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I3(\main_shift64RightJammingexit9ii_95_reg[26]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[26]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[26]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[26]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[27]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[28]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[27]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [27]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit9ii_95_reg[27]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[27]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[29]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[27]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[27]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[28]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[29]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[28]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [28]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexit9ii_95_reg[28]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[28]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[30]_i_4_n_0 ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[28]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[28]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [4]),
        .O(\main_shift64RightJammingexit9ii_95_reg[28]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[29]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[30]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[29]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [29]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[29]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[31]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[29]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_95_reg[29]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[25]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[2]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[3]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[2]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[2]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[4]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[2]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[2]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_17_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[30]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[31]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[30]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [30]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[30]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[32]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[30]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_95_reg[30]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[26]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[31]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[32]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[31]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [31]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[31]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[33]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[31]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_95_reg[31]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[27]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[32]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[33]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[32]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [32]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[32]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[34]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[32]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexit9ii_95_reg[32]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I1(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[28]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[33]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[34]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[33]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [33]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[33]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[35]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[33]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[33]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[33]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[34]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[35]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[34]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [34]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[34]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[36]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[34]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[34]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[34]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[35]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[36]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[35]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [35]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[35]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[37]_i_5_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[35]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[35]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[35]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[36]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[37]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[36]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [36]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[36]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[38]_i_5_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[36]_i_4_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexit9ii_95_reg[36]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [3]),
        .O(\main_shift64RightJammingexit9ii_95_reg[36]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[37]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[38]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[37]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [37]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[37]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[37]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[37]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_95_reg[37]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_95_reg[37]_i_5 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[37]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[38]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[39]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[38]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [38]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexit9ii_95_reg[38]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[38]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [1]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[38]_i_5_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_95_reg[38]_i_4 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexit9ii_95_reg[38]_i_5 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [2]),
        .O(\main_shift64RightJammingexit9ii_95_reg[38]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[39]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_8_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[39]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [39]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit9ii_95_reg[39]_i_3 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[3]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[4]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[3]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[3]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[5]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[3]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[3]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_13_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF2)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_4_n_0 ),
        .I1(\main_normalizeRoundAndPackFloat64exitii_shiftCount1iiiii_reg[4]_i_2_n_0 ),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit9ii_94_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_10 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(main_158_160_reg),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_12 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h20202F20)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_8_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I3(\main_inst/main_15_19_reg [40]),
        .I4(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_inst/main_shift64RightJammingexit9ii_95 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001000)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_5 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .I1(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0200000000000000)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_12_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_8 
       (.I0(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000002)) 
    \main_shift64RightJammingexit9ii_95_reg[40]_i_9 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(main_float64_addexit_220_reg),
        .O(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[4]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[5]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[4]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[4]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[4]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[4]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_18_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[5]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[6]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[5]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[5]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[5]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[5]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_14_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[6]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[7]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[6]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[6]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[6]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_16_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[7]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[7]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[7]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexit9ii_95_reg[7]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_12_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I5(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_1 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_2_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_10 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_18_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_11 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_19_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_12 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_13 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_14 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_15 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[9] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_16 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[14] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_17 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_ ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_18 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_19 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I3(\main_inst/main_27_30_reg_reg_n_0_[40] ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_3 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [2]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[8]_i_10_n_0 ),
        .I4(\main_shift64RightJammingexit9ii_95_reg[8]_i_11_n_0 ),
        .I5(\main_inst/main_27_expDiff0i2i_reg [1]),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_4 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_12_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_5 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_13_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_6 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_14_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_7 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_15_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_8 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_16_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexit9ii_95_reg[8]_i_9 
       (.I0(\main_inst/main_27_30_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [4]),
        .I2(\main_inst/main_27_30_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_27_expDiff0i2i_reg [5]),
        .I4(\main_inst/main_27_expDiff0i2i_reg [3]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[8]_i_17_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[8]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800B8FFB800)) 
    \main_shift64RightJammingexit9ii_95_reg[9]_i_2 
       (.I0(\main_shift64RightJammingexit9ii_95_reg[10]_i_3_n_0 ),
        .I1(\main_inst/main_27_expDiff0i2i_reg [0]),
        .I2(\main_shift64RightJammingexit9ii_95_reg[8]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexit9ii_95_reg[40]_i_9_n_0 ),
        .I4(\main_inst/main_15_19_reg [9]),
        .I5(\main_shift64RightJammingexit9ii_95_reg[40]_i_10_n_0 ),
        .O(\main_shift64RightJammingexit9ii_95_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_13 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_0 ),
        .CO(main_shift64RightJammingexit9ii_95_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_31_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_32_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_33_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_34_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_36_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_37_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_38_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_39_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_1 ,\main_inst/main_45_47 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_30_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_64_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_65_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_66_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_67_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_35_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_69_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_70_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_71_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_72_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_0 ,\main_inst/main_35_43 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_9_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_10_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_68_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_115_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_116_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_117_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_118_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7 
       (.CI(main_shift64RightJammingexit9ii_95_reg_reg[3]),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_14_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_15_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8 
       (.CI(\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_17_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_0 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_1 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_2 ,\main_shift64RightJammingexit9ii_95_reg_reg[0]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexit9ii_95_reg[0]_i_18_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_19_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_20_n_0 ,\main_shift64RightJammingexit9ii_95_reg[0]_i_21_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    main_shift64RightJammingexit9ii_99_reg_i_1
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_[1] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(main_float64_addexit_220_reg),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_inst/main_shift64RightJammingexit9ii_99_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[11]_i_11 
       (.I0(\main_inst/A [7]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [7]),
        .O(main_shift64RightJammingexit9ii_ii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[11]_i_12 
       (.I0(\main_inst/A [6]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [6]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[11]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[11]_i_13 
       (.I0(\main_inst/A [5]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [5]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[11]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[11]_i_14 
       (.I0(\main_inst/A [4]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [4]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[11]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[15]_i_11 
       (.I0(\main_inst/A [11]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [11]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[15]_i_12 
       (.I0(\main_inst/A [10]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [10]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[15]_i_13 
       (.I0(\main_inst/A [9]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [9]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[15]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[15]_i_14 
       (.I0(\main_inst/A [8]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [8]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[15]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[19]_i_11 
       (.I0(\main_inst/A [15]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [15]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[19]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[19]_i_12 
       (.I0(\main_inst/A [14]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [14]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[19]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[19]_i_13 
       (.I0(\main_inst/A [13]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [13]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[19]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[19]_i_14 
       (.I0(\main_inst/A [12]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [12]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[19]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[23]_i_11 
       (.I0(\main_inst/A [19]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [19]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[23]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[23]_i_12 
       (.I0(\main_inst/A [18]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [18]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[23]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[23]_i_13 
       (.I0(\main_inst/A [17]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [17]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[23]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[23]_i_14 
       (.I0(\main_inst/A [16]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [16]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[23]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[27]_i_11 
       (.I0(\main_inst/A [23]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [23]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[27]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[27]_i_12 
       (.I0(\main_inst/A [22]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [22]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[27]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[27]_i_13 
       (.I0(\main_inst/A [21]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [21]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[27]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[27]_i_14 
       (.I0(\main_inst/A [20]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [20]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[27]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[31]_i_11 
       (.I0(\main_inst/A [27]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [27]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[31]_i_12 
       (.I0(\main_inst/A [26]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [26]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[31]_i_13 
       (.I0(\main_inst/A [25]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [25]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[31]_i_14 
       (.I0(\main_inst/A [24]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [24]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[35]_i_11 
       (.I0(\main_inst/A [31]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [31]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[35]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[35]_i_12 
       (.I0(\main_inst/A [30]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [30]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[35]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[35]_i_13 
       (.I0(\main_inst/A [29]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [29]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[35]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[35]_i_14 
       (.I0(\main_inst/A [28]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [28]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[35]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[39]_i_11 
       (.I0(\main_inst/A [35]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [35]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[39]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[39]_i_12 
       (.I0(\main_inst/A [34]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [34]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[39]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[39]_i_13 
       (.I0(\main_inst/A [33]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [33]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[39]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[39]_i_14 
       (.I0(\main_inst/A [32]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [32]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[39]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[43]_i_10 
       (.I0(\main_inst/A [37]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [37]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[43]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[43]_i_11 
       (.I0(\main_inst/A [36]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [36]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[43]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[43]_i_8 
       (.I0(\main_inst/A [39]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [39]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[43]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[43]_i_9 
       (.I0(\main_inst/A [38]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [38]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[43]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[48]_i_5 
       (.I0(\main_inst/A [40]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [40]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[48]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[7]_i_11 
       (.I0(\main_inst/A [3]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [3]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[7]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[7]_i_12 
       (.I0(\main_inst/A [2]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [2]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[7]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[7]_i_13 
       (.I0(\main_inst/A [1]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [1]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[7]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \main_shift64RightJammingexit9ii_ii_reg[7]_i_14 
       (.I0(\main_inst/A [0]),
        .I1(\main_inst/main_shift64RightJammingexit9ii_95_reg [0]),
        .O(\main_shift64RightJammingexit9ii_ii_reg[7]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_178,ZERO_177,ZERO_176,ZERO_175}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_7 }),
        .S(\main_inst/C [11:8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_0 ),
        .CO(main_shift64RightJammingexit9ii_ii_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [7:4]),
        .O(\main_inst/C [8:5]),
        .S({main_shift64RightJammingexit9ii_ii_reg,\main_shift64RightJammingexit9ii_ii_reg[11]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[11]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[11]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[11]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_174,ZERO_173,ZERO_172,ZERO_171}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_7 }),
        .S(\main_inst/C [15:12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10 
       (.CI(main_shift64RightJammingexit9ii_ii_reg_reg[3]),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [11:8]),
        .O(\main_inst/C [12:9]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[15]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[15]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[15]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[15]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_170,ZERO_169,ZERO_168,ZERO_167}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_7 }),
        .S(\main_inst/C [19:16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[15]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [15:12]),
        .O(\main_inst/C [16:13]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[19]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[19]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[19]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[19]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_166,ZERO_165,ZERO_164,ZERO_163}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_7 }),
        .S(\main_inst/C [23:20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[19]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [19:16]),
        .O(\main_inst/C [20:17]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[23]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[23]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[23]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[23]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_162,ZERO_161,ZERO_160,ZERO_159}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_7 }),
        .S(\main_inst/C [27:24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[23]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [23:20]),
        .O(\main_inst/C [24:21]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[27]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[27]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[27]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[27]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_158,ZERO_157,ZERO_156,ZERO_155}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_7 }),
        .S(\main_inst/C [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[27]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [27:24]),
        .O(\main_inst/C [28:25]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[31]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[31]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[31]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[31]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_154,ZERO_153,ZERO_152,ZERO_151}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_7 }),
        .S(\main_inst/C [35:32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[31]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [31:28]),
        .O(\main_inst/C [32:29]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[35]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[35]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[35]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[35]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_150,ZERO_149,ZERO_148,ZERO_147}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_7 }),
        .S(\main_inst/C [39:36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[35]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [35:32]),
        .O(\main_inst/C [36:33]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[39]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[39]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[39]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[39]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_146,ZERO_145,ZERO_144,ZERO_143}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_7 }),
        .S({\main_inst/C [3:1],ZERO_136}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,ZERO_142}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_1_n_7 }),
        .S({ZERO_249,\main_inst/C [42:40]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[39]_i_10_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [39:36]),
        .O(\main_inst/C [40:37]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[43]_i_8_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[43]_i_9_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[43]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[43]_i_11_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[48]_i_4 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[43]_i_7_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/A [40]}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[48]_i_4_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[48]_i_4_n_5 ,\main_inst/C [42:41]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\main_shift64RightJammingexit9ii_ii_reg[48]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC \main_shift64RightJammingexit9ii_ii_reg_reg[63]_i_1_VCC 
       (.P(\main_shift64RightJammingexit9ii_ii_reg_reg[63]_i_1_VCC_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1 
       (.CI(\main_shift64RightJammingexit9ii_ii_reg_reg[3]_i_1_n_0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({ZERO_140,ZERO_139,ZERO_138,ZERO_137}),
        .O({\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_4 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_5 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_6 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_1_n_7 }),
        .S(\main_inst/C [7:4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_0 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_1 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_2 ,\main_shift64RightJammingexit9ii_ii_reg_reg[7]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI(\main_inst/A [3:0]),
        .O(\main_inst/C [4:1]),
        .S({\main_shift64RightJammingexit9ii_ii_reg[7]_i_11_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[7]_i_12_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[7]_i_13_n_0 ,\main_shift64RightJammingexit9ii_ii_reg[7]_i_14_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_10 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_7_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_100 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(main_shift64RightJammingexitii_z0iii_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_101 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_102 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_155_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_103 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_156_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_104 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_105 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_107 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_108 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_109 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_110 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_111 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_161_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_126_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_162_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_163_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_111_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_112 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_164_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_163_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_165_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_166_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000050300010F01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_113 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_167_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_166_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_168_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_169_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3FFFFFFCFFFFFFFD)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_114 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_170_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .I4(\main_inst/main_169_expDiff1ii_reg [0]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_171_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_115 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_172_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_116 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_173_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_117 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_172_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_118 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_173_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_119 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_176_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_119_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h400143C17C3D7FFD))
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_120 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_177_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_120_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_121 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_178_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_176_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_121_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_122 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_179_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_177_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_122_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_123 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_178_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_180_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_123_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_124 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_179_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_181_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_124_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_125 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_180_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_182_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_125_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_126 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_181_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_183_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_126_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_127 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_85_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_184_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_127_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_128 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_149_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_185_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_128_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_129 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_186_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_129_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_13 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_31_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_24_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_32_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_33_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_130 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_187_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_131 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_188_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_132 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_184_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_189_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_132_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_133 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_185_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_190_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_133_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_134 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_135 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_136 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_189_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_191_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_136_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_137 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_190_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_192_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_137_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_138 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_139 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_14 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_34_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_33_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_35_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_36_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_140 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_193_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_140_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_141 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_194_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_142 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_143 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_144 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_145 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_195_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_145_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_146 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_196_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_146_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_147 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_147_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_148 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_148_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_149 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_197_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_149_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_15 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_37_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_36_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_38_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_39_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_150 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_150_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_151 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_151_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_152 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_152_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_153 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_153_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_154 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_154_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_155 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_155_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_156 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_156_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_157 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_157_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_158 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_158_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_159 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_159_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_16 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_40_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_39_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_41_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_42_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_160 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_160_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_161 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_182_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_198_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_161_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_162 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_183_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_199_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_162_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_163 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_198_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_200_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_163_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_164 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_199_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_201_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_164_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBE82828282828282)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_165 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_200_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_202_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_165_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBE82828282828282)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_166 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_201_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_203_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_166_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_167 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_167_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBC80000000000202)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_168 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_203_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_171_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_168_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_169 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_169_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFE2B80000E2)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_17 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_43_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_44_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_inst/main_169_expDiff1ii_reg [1]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_45_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_170 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_170_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_171 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_171_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_172 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_191_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_205_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_172_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_173 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_192_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_206_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_173_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_174 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_174_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_175 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_175_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_176 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_205_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_207_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_176_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_177 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_206_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_208_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_177_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_178 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_178_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_179 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_179_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFFFE2B80000E2)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_18 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_46_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_47_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_inst/main_169_expDiff1ii_reg [1]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_48_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_180 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_207_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_180_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_181 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_208_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_181_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_182 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_178_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_182_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB888888888888888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_183 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_179_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_183_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_184 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_209_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_184_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_185 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_210_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_185_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_186 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_186_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_187 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_187_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_188 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_188_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_189 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_189_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_19 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_44_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_45_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_190 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_190_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_191 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_191_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFC00000A0C00000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_192 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_192_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_193 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_193_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_194 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_194_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_195 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_195_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_196 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_196_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_197 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_197_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_198 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_198_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_199 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_199_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEAEFFFFFEAE0000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_2 
       (.I0(\main_inst/main_177_185 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_4_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[1]_i_2_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I5(\main_inst/main_187_189 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_20 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_47_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_48_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_200 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_200_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB000800000000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_201 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_201_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_202 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_202_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h80)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_203 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_203_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_204 
       (.I0(\main_inst/main_169_expDiff1ii_reg [1]),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [2]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_204_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0008000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_205 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_205_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0008000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_206 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_206_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_207 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_207_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB0800000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_208 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_208_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_209 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_209_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_21 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_44_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_51_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_210 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_210_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_22 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_47_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_52_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_23 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_53_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_51_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_24 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_52_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_27 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_64_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_42_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_65_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_66_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_28 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_67_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_66_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_68_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_69_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_29 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_70_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_69_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_71_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_72_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_30 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_73_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_72_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_74_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_75_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_31 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_53_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_76_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_32 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_77_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_33 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_76_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_78_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_34 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_77_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_35 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_80_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_78_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_36 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_82_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_37 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_80_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_83_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_38 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_82_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_39 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_85_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_83_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_4 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[2]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[4]_i_3_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_10_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_40 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_86_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_41 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_85_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_87_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_42 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_86_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_43 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_92_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_44 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_93_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_45 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_94_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_95_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_46 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_96_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_47 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_97_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_48 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_98_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_99_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_49 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(main_shift64RightJammingexitii_z0iii_reg),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_50 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_101_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_51 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_95_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_102_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_52 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_99_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_103_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_53 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_104_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_54 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_105_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_56 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_57 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_58 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_60 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_115_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_75_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_116_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_117_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_61 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_118_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_117_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_119_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_120_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_62 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_121_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_120_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_122_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_123_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_63 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_124_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_123_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_125_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_126_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hBE82)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_64 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_87_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_127_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_65 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_128_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_66 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_129_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_127_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_67 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_128_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_68 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_129_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_132_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_68_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_69 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_133_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_7 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_17_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_18_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_70 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_132_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_71 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_133_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_72 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_130_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_136_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBFFEBC3E83C28002)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_73 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_131_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_137_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_73_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_74 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_134_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_138_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_136_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEBFFEBC3283C2800)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_75 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_135_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_139_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_137_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_76 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_102_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_80_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_77 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_103_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_140_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_78 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_53_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_141_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_79 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_142_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_8 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_19_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_18_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_20_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_21_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_80 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_143_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_81 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_144_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_82 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_140_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_145_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_83 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_141_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_146_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3088FFFF30880000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_84 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_147_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_85 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_148_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_86 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_145_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_149_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hABFEA802)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_87 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_146_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_129_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_88 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_150_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFE0001)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_89 
       (.I0(\main_inst/main_169_expDiff1ii_reg [3]),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [2]),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010501)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_9 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[0]_i_22_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_21_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_23_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [0]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_24_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFE00000001)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_90 
       (.I0(\main_inst/main_169_expDiff1ii_reg [4]),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_inst/main_169_expDiff1ii_reg [1]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_91 
       (.I0(\main_inst/main_169_expDiff1ii_reg [2]),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_92 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_93 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_94 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_151_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_95 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_152_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_96 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_97 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_98 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_153_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h3808FFFF38080000)) 
    \main_shift64RightJammingexitii_z0iii_reg[0]_i_99 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[0]_i_89_n_0 ),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[0]_i_90_n_0 ),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[0]_i_91_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[0]_i_154_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[0]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[10]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[10]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[11]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[10]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[12]_i_3_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [1]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[8]_i_2_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[11]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[11]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[12]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[11]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[11]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[11]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[11]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[11] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[12]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[12]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[13]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[12]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[14]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[12]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[12]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[12]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[12]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[12] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[13]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[13]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[14]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[13]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[13]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[13]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[13]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[13] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[14]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[14]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[15]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[14]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[14]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[14]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[14]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[14]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[14] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[15]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[15]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[16]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[15]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[15]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[15]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[15]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[15] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[16]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[16]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[17]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[16]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[16]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[16]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[16]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[17]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[17]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[18]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[17]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[17]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[17]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[17]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[18]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[18]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[19]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[18]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[18]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[19]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[19]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[20]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[19]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[19]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[1]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[2]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[1]_i_2_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [0]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8FFB833B8CCB800)) 
    \main_shift64RightJammingexitii_z0iii_reg[1]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[3]_i_3_n_0 ),
        .I3(\main_inst/main_169_expDiff1ii_reg [1]),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[5]_i_3_n_0 ),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[1]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[1]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[9]_i_15_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[20]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[20]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[21]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[20]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[20]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[21]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[21]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[22]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[21]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[21]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[22]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[22]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[23]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[22]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[22]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[23]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[23]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[24]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[23]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[23]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[24]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[24]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[25]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[24]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[26]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[24]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[25]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[25]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[26]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[25]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[27]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \main_shift64RightJammingexitii_z0iii_reg[25]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I5(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[26]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[26]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[27]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[26]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[28]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[26]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[26]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[30] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[26]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[27]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[27]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[28]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \main_shift64RightJammingexitii_z0iii_reg[27]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[29]_i_3_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [1]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[27]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[27]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[31] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[27]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[27] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[28]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[28]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[29]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[28]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[28]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[30]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[28]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[28]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[28] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[29]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[29]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[30]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[29]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[29]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[31]_i_3_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[29]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[29]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[29] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [4]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexitii_z0iii_reg[2]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[2]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [0]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[3]_i_2_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[2]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[6]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[2]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[2]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_6_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[30]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[30]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[31]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[30]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[32]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[30]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexitii_z0iii_reg[30]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [4]),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[26]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[31]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[31]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[32]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[31]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[33]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[31]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexitii_z0iii_reg[31]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [4]),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[27]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[32]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[32]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[33]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[32]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[34]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[32]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexitii_z0iii_reg[32]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [4]),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[28]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[33]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[33]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[34]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[33]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[35]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[33]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \main_shift64RightJammingexitii_z0iii_reg[33]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [4]),
        .I1(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_expDiff1ii_reg [3]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[29]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[34]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[34]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[35]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[34]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[36]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[34]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[34]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [4]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[35]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[35]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[36]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[35]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[37]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[35]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[35]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [4]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[36]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[36]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[37]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[36]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[38]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[36]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[36]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [4]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[37]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[37]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[38]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[37]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[39]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[37]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \main_shift64RightJammingexitii_z0iii_reg[37]_i_3 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_inst/main_169_expDiff1ii_reg [4]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_expDiff1ii_reg [3]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[38]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[38]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[39]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[38]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[38]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[38]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[38]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [3]),
        .I1(\main_inst/main_169_expDiff1ii_reg [5]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[38]_i_4 
       (.I0(\main_inst/main_169_expDiff1ii_reg [3]),
        .I1(\main_inst/main_169_expDiff1ii_reg [5]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[39]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[39]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[40]_i_2_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[39]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[39]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[39]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[39]_i_3 
       (.I0(\main_inst/main_169_expDiff1ii_reg [3]),
        .I1(\main_inst/main_169_expDiff1ii_reg [5]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[39]_i_4 
       (.I0(\main_inst/main_169_expDiff1ii_reg [3]),
        .I1(\main_inst/main_169_expDiff1ii_reg [5]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [2]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[3]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[3]_i_2_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [0]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[3]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[5]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[3]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[3]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[11]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[19] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[35] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[40]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[40]_i_2_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_5_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[40]_i_2 
       (.I0(\main_inst/main_169_expDiff1ii_reg [2]),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0048)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[41]_i_3_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [0]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[41]_i_5_n_0 ),
        .O(\main_inst/main_shift64RightJammingexitii_z0iii [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0004)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000400)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_5 
       (.I0(\main_inst/main_169_expDiff1ii_reg [2]),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[41]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \main_shift64RightJammingexitii_z0iii_reg[41]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[6] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[41]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexitii_z0iii_reg[4]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [0]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[5]_i_2_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[4]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_5_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[4]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[4]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[12]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[20] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[36] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[5]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[5]_i_2_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [0]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[5]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[5]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[5]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[13]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[21] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[37] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexitii_z0iii_reg[6]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [0]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[7]_i_2_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[6]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[6]_i_3_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[6]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[14]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[22] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[38] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800B800FF000000)) 
    \main_shift64RightJammingexitii_z0iii_reg[7]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[7]_i_2_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [0]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[7]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h88BBB8888888B888)) 
    \main_shift64RightJammingexitii_z0iii_reg[7]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[15]_i_4_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [3]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[23] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [4]),
        .I4(\main_inst/main_169_expDiff1ii_reg [5]),
        .I5(\main_inst/main_169_172_reg_reg_n_0_[39] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF00B8000000B800)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_1 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[8]_i_2_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [1]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I4(\main_inst/main_169_expDiff1ii_reg [0]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[9]_i_5_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[14]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[8]_i_4_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_3 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[12]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[8]_i_5_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_4 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[34] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[18] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[8]_i_6_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_5 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[32] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[16] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[8]_i_7_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_6 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[26] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_ ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[8]_i_7 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[24] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[40] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[8]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \main_shift64RightJammingexitii_z0iii_reg[9]_i_10 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[33] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_172_reg_reg_n_0_[17] ),
        .I3(\main_inst/main_169_expDiff1ii_reg [5]),
        .I4(\main_inst/main_169_expDiff1ii_reg [3]),
        .I5(\main_shift64RightJammingexitii_z0iii_reg[9]_i_15_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3808)) 
    \main_shift64RightJammingexitii_z0iii_reg[9]_i_15 
       (.I0(\main_inst/main_169_172_reg_reg_n_0_[25] ),
        .I1(\main_inst/main_169_expDiff1ii_reg [4]),
        .I2(\main_inst/main_169_expDiff1ii_reg [5]),
        .I3(\main_inst/main_169_172_reg_reg_n_0_[41] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[9]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hA808)) 
    \main_shift64RightJammingexitii_z0iii_reg[9]_i_2 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[41]_i_4_n_0 ),
        .I1(\main_shift64RightJammingexitii_z0iii_reg[9]_i_5_n_0 ),
        .I2(\main_inst/main_169_expDiff1ii_reg [0]),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[10]_i_2_n_0 ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h20)) 
    \main_shift64RightJammingexitii_z0iii_reg[9]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .O(\main_shift64RightJammingexitii_z0iii_reg[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \main_shift64RightJammingexitii_z0iii_reg[9]_i_5 
       (.I0(\main_shift64RightJammingexitii_z0iii_reg[15]_i_3_n_0 ),
        .I1(\main_inst/main_169_expDiff1ii_reg [2]),
        .I2(\main_shift64RightJammingexitii_z0iii_reg[11]_i_3_n_0 ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[13]_i_3_n_0 ),
        .I4(\main_shift64RightJammingexitii_z0iii_reg[9]_i_10_n_0 ),
        .I5(\main_inst/main_169_expDiff1ii_reg [1]),
        .O(\main_shift64RightJammingexitii_z0iii_reg[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_106 
       (.CI(\<const0>__0__0 ),
        .CO(main_shift64RightJammingexitii_z0iii_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_157_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_158_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_159_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_160_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_27_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_28_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_29_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_30_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_25_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const1>__0__0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_56_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_57_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_58_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_26_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_60_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_61_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_62_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_63_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_0 ,\main_inst/main_177_185 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_7_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_8_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_9_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_11_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_1 ,\main_inst/main_187_189 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55 
       (.CI(main_shift64RightJammingexitii_z0iii_reg_reg[3]),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_55_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_107_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_108_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_109_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_110_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59 
       (.CI(\<const0>__0__0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_59_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_111_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_112_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_113_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_114_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6 
       (.CI(\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_12_n_0 ),
        .CO({\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_0 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_1 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_2 ,\main_shift64RightJammingexitii_z0iii_reg_reg[0]_i_6_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\main_shift64RightJammingexitii_z0iii_reg[0]_i_13_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_14_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_15_n_0 ,\main_shift64RightJammingexitii_z0iii_reg[0]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000010055550100)) 
    memory_controller_enable_reg_a_i_1
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg ),
        .I3(memory_controller_enable_reg_a_i_2_n_0),
        .I4(\main_inst/cur_state_reg_n_0_ ),
        .I5(memory_controller_enable_reg_a_i_3_n_0),
        .O(memory_controller_enable_a));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    memory_controller_enable_reg_a_i_2
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .O(memory_controller_enable_reg_a_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEEEFEFBF7EFF7E)) 
    memory_controller_enable_reg_a_i_3
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg ),
        .I4(\main_inst/roundAndPackFloat64_memory_controller_enable_a ),
        .I5(\main_inst/cur_state_reg_n_0_[5] ),
        .O(memory_controller_enable_reg_a_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001C54)) 
    memory_controller_enable_reg_a_i_4
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_enable_a ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000200000000)) 
    memory_controller_enable_reg_b_i_1
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(memory_controller_enable_reg_b_i_2_n_0),
        .O(memory_controller_enable_b));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1811)) 
    memory_controller_enable_reg_b_i_2
       (.I0(\main_inst/cur_state_reg ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .O(memory_controller_enable_reg_b_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* CLOCK_DOMAINS = "COMMON" *) 
  (* IS_CLOCK_GATED *) 
  (* METHODOLOGY_DRC_VIOS = "{SYNTH-6 {cell *THIS*}} {SYNTH-7 {cell *THIS*}}" *) 
  (* POWER_OPTED_CE = "ENBWREN=NEW" *) 
  (* RTL_RAM_BITS = "32" *) 
  (* RTL_RAM_NAME = "ram" *) 
  (* bram_addr_begin = "0" *) 
  (* bram_addr_end = "1023" *) 
  (* bram_slice_begin = "0" *) 
  (* bram_slice_end = "35" *) 
  RAMB36E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .EN_ECC_READ("FALSE"),
    .EN_ECC_WRITE("FALSE"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_40(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_41(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_42(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_43(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_44(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_45(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_46(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_47(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_48(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_49(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_4F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_50(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_51(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_52(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_53(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_54(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_55(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_56(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_57(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_58(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_59(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_5F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_60(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_61(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_62(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_63(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_64(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_65(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_66(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_67(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_68(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_69(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_6F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_70(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_71(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_72(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_73(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_74(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_75(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_76(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_77(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_78(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_79(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_7F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_A(36'h000000000),
    .INIT_B(36'h000000000),
    .INIT_FILE("NONE"),
    .IS_CLKARDCLK_INVERTED(1'b0),
    .IS_CLKBWRCLK_INVERTED(1'b0),
    .IS_ENARDEN_INVERTED(1'b0),
    .IS_ENBWREN_INVERTED(1'b0),
    .IS_RSTRAMARSTRAM_INVERTED(1'b0),
    .IS_RSTRAMB_INVERTED(1'b0),
    .IS_RSTREGARSTREG_INVERTED(1'b0),
    .IS_RSTREGB_INVERTED(1'b0),
    .RAM_EXTENSION_A("NONE"),
    .RAM_EXTENSION_B("NONE"),
    .RAM_MODE("TDP"),
    .RDADDR_COLLISION_HWCONFIG("DELAYED_WRITE"),
    .READ_WIDTH_A(36),
    .READ_WIDTH_B(36),
    .RSTREG_PRIORITY_A("RSTREG"),
    .RSTREG_PRIORITY_B("RSTREG"),
    .SIM_COLLISION_CHECK("ALL"),
    .SIM_DEVICE("7SERIES"),
    .SRVAL_A(36'h000000000),
    .SRVAL_B(36'h000000000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(36),
    .WRITE_WIDTH_B(36)) 
    \memory_controller_inst/float_exception_flags/ram_reg 
       (.ADDRARDADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .ADDRBWRADDR({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .CASCADEINA(\<const1>__0__0 ),
        .CASCADEINB(\<const1>__0__0 ),
        .CLKARDCLK(clk),
        .CLKBWRCLK(clk),
        .DIADI({ram_reg_i_1_n_0,ram_reg_i_2_n_0,ram_reg_i_3_n_0,ram_reg_i_4_n_0,ram_reg_i_5_n_0,ram_reg_i_6_n_0,ram_reg_i_7_n_0,ram_reg_i_8_n_0,ram_reg_i_9_n_0,ram_reg_i_10_n_0,ram_reg_i_11_n_0,ram_reg_i_12_n_0,ram_reg_i_13_n_0,ram_reg_i_14_n_0,ram_reg_i_15_n_0,ram_reg_i_16_n_0,ram_reg_i_17_n_0,ram_reg_i_18_n_0,ram_reg_i_19_n_0,ram_reg_i_20_n_0,ram_reg_i_21_n_0,ram_reg_i_22_n_0,ram_reg_i_23_n_0,ram_reg_i_24_n_0,ram_reg_i_25_n_0,ram_reg_i_26_n_0,ram_reg_i_27_n_0,memory_controller_in_a,ram_reg_i_29_n_0,ram_reg_i_30_n_0,ram_reg_i_31_n_0,ram_reg_i_32_n_0}),
        .DIBDI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPADIP({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .DIPBDIP({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .DOADO(\memory_controller_inst/float_exception_flags/q_a_wire ),
        .DOBDO(\memory_controller_inst/float_exception_flags/q_b_wire ),
        .ENARDEN(\<const1>__0__0 ),
        .ENBWREN(\memory_controller_inst/float_exception_flags/ram_reg_ENBWREN_cooolgate_en_sig_1 ),
        .REGCEAREGCE(\<const0>__0__0 ),
        .REGCEB(\<const0>__0__0 ),
        .RSTRAMARSTRAM(\<const0>__0__0 ),
        .RSTRAMB(\<const0>__0__0 ),
        .RSTREGARSTREG(\<const0>__0__0 ),
        .RSTREGB(\<const0>__0__0 ),
        .WEA({\memory_controller_inst/float_exception_flags_write_enable_a ,\memory_controller_inst/float_exception_flags_write_enable_a ,\memory_controller_inst/float_exception_flags_write_enable_a ,\memory_controller_inst/float_exception_flags_write_enable_a }),
        .WEBWE({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \memory_controller_inst/float_exception_flags/ram_reg_ENBWREN_cooolgate_en_gate_1 
       (.I0(\select_float_exception_flags_reg_b[1]_i_5_n_0 ),
        .I1(\select_float_exception_flags_reg_b[1]_i_3_n_0 ),
        .I2(memory_controller_address_b),
        .O(\memory_controller_inst/float_exception_flags/ram_reg_ENBWREN_cooolgate_en_sig_1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_enable_reg_a_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(memory_controller_enable_a),
        .Q(\memory_controller_inst/memory_controller_enable_reg_a ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_enable_reg_b_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(memory_controller_enable_b),
        .Q(\memory_controller_inst/memory_controller_enable_reg_b ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [0]),
        .Q(memory_controller_out_a[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [10]),
        .Q(memory_controller_out_a[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [11]),
        .Q(memory_controller_out_a[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [12]),
        .Q(memory_controller_out_a[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [13]),
        .Q(memory_controller_out_a[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [14]),
        .Q(memory_controller_out_a[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [15]),
        .Q(memory_controller_out_a[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [16]),
        .Q(memory_controller_out_a[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [17]),
        .Q(memory_controller_out_a[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [18]),
        .Q(memory_controller_out_a[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [19]),
        .Q(memory_controller_out_a[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [1]),
        .Q(memory_controller_out_a[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [20]),
        .Q(memory_controller_out_a[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [21]),
        .Q(memory_controller_out_a[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [22]),
        .Q(memory_controller_out_a[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [23]),
        .Q(memory_controller_out_a[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [24]),
        .Q(memory_controller_out_a[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [25]),
        .Q(memory_controller_out_a[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [26]),
        .Q(memory_controller_out_a[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [27]),
        .Q(memory_controller_out_a[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [28]),
        .Q(memory_controller_out_a[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [29]),
        .Q(memory_controller_out_a[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [2]),
        .Q(memory_controller_out_a[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [30]),
        .Q(memory_controller_out_a[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [31]),
        .Q(memory_controller_out_a[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [3]),
        .Q(memory_controller_out_a[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [4]),
        .Q(memory_controller_out_a[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [5]),
        .Q(memory_controller_out_a[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [6]),
        .Q(memory_controller_out_a[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [7]),
        .Q(memory_controller_out_a[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [8]),
        .Q(memory_controller_out_a[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_a_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_a [9]),
        .Q(memory_controller_out_a[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [0]),
        .Q(memory_controller_out_b[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [10]),
        .Q(memory_controller_out_b[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [11]),
        .Q(memory_controller_out_b[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[12] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [12]),
        .Q(memory_controller_out_b[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[13] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [13]),
        .Q(memory_controller_out_b[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[14] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [14]),
        .Q(memory_controller_out_b[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[15] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [15]),
        .Q(memory_controller_out_b[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[16] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [16]),
        .Q(memory_controller_out_b[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[17] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [17]),
        .Q(memory_controller_out_b[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[18] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [18]),
        .Q(memory_controller_out_b[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[19] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [19]),
        .Q(memory_controller_out_b[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [1]),
        .Q(memory_controller_out_b[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[20] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [20]),
        .Q(memory_controller_out_b[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[21] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [21]),
        .Q(memory_controller_out_b[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[22] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [22]),
        .Q(memory_controller_out_b[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[23] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [23]),
        .Q(memory_controller_out_b[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[24] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [24]),
        .Q(memory_controller_out_b[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[25] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [25]),
        .Q(memory_controller_out_b[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[26] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [26]),
        .Q(memory_controller_out_b[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[27] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [27]),
        .Q(memory_controller_out_b[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[28] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [28]),
        .Q(memory_controller_out_b[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[29] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [29]),
        .Q(memory_controller_out_b[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [2]),
        .Q(memory_controller_out_b[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[30] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [30]),
        .Q(memory_controller_out_b[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[31] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [31]),
        .Q(memory_controller_out_b[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [3]),
        .Q(memory_controller_out_b[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [4]),
        .Q(memory_controller_out_b[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [5]),
        .Q(memory_controller_out_b[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [6]),
        .Q(memory_controller_out_b[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [7]),
        .Q(memory_controller_out_b[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [8]),
        .Q(memory_controller_out_b[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/memory_controller_out_reg_b_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\memory_controller_inst/memory_controller_out_b [9]),
        .Q(memory_controller_out_b[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/select_float_exception_flags_reg_a_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\select_float_exception_flags_reg_a[1]_i_1_n_0 ),
        .Q(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \memory_controller_inst/select_float_exception_flags_reg_b_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\select_float_exception_flags_reg_b[1]_i_1_n_0 ),
        .Q(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[0]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [0]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[0]),
        .O(\memory_controller_inst/memory_controller_out_a [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[10]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [10]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[10]),
        .O(\memory_controller_inst/memory_controller_out_a [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[11]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [11]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[11]),
        .O(\memory_controller_inst/memory_controller_out_a [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[12]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [12]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[12]),
        .O(\memory_controller_inst/memory_controller_out_a [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[13]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [13]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[13]),
        .O(\memory_controller_inst/memory_controller_out_a [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[14]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [14]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[14]),
        .O(\memory_controller_inst/memory_controller_out_a [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[15]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [15]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[15]),
        .O(\memory_controller_inst/memory_controller_out_a [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[16]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [16]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[16]),
        .O(\memory_controller_inst/memory_controller_out_a [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[17]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [17]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[17]),
        .O(\memory_controller_inst/memory_controller_out_a [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[18]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [18]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[18]),
        .O(\memory_controller_inst/memory_controller_out_a [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[19]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [19]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[19]),
        .O(\memory_controller_inst/memory_controller_out_a [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[1]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [1]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[1]),
        .O(\memory_controller_inst/memory_controller_out_a [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[20]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [20]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[20]),
        .O(\memory_controller_inst/memory_controller_out_a [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[21]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [21]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[21]),
        .O(\memory_controller_inst/memory_controller_out_a [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[22]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [22]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[22]),
        .O(\memory_controller_inst/memory_controller_out_a [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[23]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [23]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[23]),
        .O(\memory_controller_inst/memory_controller_out_a [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[24]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [24]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[24]),
        .O(\memory_controller_inst/memory_controller_out_a [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[25]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [25]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[25]),
        .O(\memory_controller_inst/memory_controller_out_a [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[26]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [26]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[26]),
        .O(\memory_controller_inst/memory_controller_out_a [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[27]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [27]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[27]),
        .O(\memory_controller_inst/memory_controller_out_a [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[28]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [28]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[28]),
        .O(\memory_controller_inst/memory_controller_out_a [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[29]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [29]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[29]),
        .O(\memory_controller_inst/memory_controller_out_a [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[2]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [2]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[2]),
        .O(\memory_controller_inst/memory_controller_out_a [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[30]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [30]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[30]),
        .O(\memory_controller_inst/memory_controller_out_a [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[31]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [31]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[31]),
        .O(\memory_controller_inst/memory_controller_out_a [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[3]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [3]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[3]),
        .O(\memory_controller_inst/memory_controller_out_a [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[4]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [4]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[4]),
        .O(\memory_controller_inst/memory_controller_out_a [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[5]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [5]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[5]),
        .O(\memory_controller_inst/memory_controller_out_a [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[6]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [6]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[6]),
        .O(\memory_controller_inst/memory_controller_out_a [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[7]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [7]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[7]),
        .O(\memory_controller_inst/memory_controller_out_a [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[8]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [8]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[8]),
        .O(\memory_controller_inst/memory_controller_out_a [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_a[9]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_a_wire [9]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_a ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_a ),
        .I3(memory_controller_out_a[9]),
        .O(\memory_controller_inst/memory_controller_out_a [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[0]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [0]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[0]),
        .O(\memory_controller_inst/memory_controller_out_b [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[10]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [10]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[10]),
        .O(\memory_controller_inst/memory_controller_out_b [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[11]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [11]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[11]),
        .O(\memory_controller_inst/memory_controller_out_b [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[12]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [12]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[12]),
        .O(\memory_controller_inst/memory_controller_out_b [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[13]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [13]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[13]),
        .O(\memory_controller_inst/memory_controller_out_b [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[14]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [14]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[14]),
        .O(\memory_controller_inst/memory_controller_out_b [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[15]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [15]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[15]),
        .O(\memory_controller_inst/memory_controller_out_b [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[16]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [16]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[16]),
        .O(\memory_controller_inst/memory_controller_out_b [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[17]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [17]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[17]),
        .O(\memory_controller_inst/memory_controller_out_b [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[18]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [18]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[18]),
        .O(\memory_controller_inst/memory_controller_out_b [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[19]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [19]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[19]),
        .O(\memory_controller_inst/memory_controller_out_b [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[1]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [1]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[1]),
        .O(\memory_controller_inst/memory_controller_out_b [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[20]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [20]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[20]),
        .O(\memory_controller_inst/memory_controller_out_b [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[21]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [21]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[21]),
        .O(\memory_controller_inst/memory_controller_out_b [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[22]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [22]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[22]),
        .O(\memory_controller_inst/memory_controller_out_b [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[23]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [23]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[23]),
        .O(\memory_controller_inst/memory_controller_out_b [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[24]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [24]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[24]),
        .O(\memory_controller_inst/memory_controller_out_b [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[25]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [25]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[25]),
        .O(\memory_controller_inst/memory_controller_out_b [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[26]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [26]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[26]),
        .O(\memory_controller_inst/memory_controller_out_b [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[27]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [27]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[27]),
        .O(\memory_controller_inst/memory_controller_out_b [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[28]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [28]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[28]),
        .O(\memory_controller_inst/memory_controller_out_b [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[29]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [29]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[29]),
        .O(\memory_controller_inst/memory_controller_out_b [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[2]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [2]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[2]),
        .O(\memory_controller_inst/memory_controller_out_b [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[30]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [30]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[30]),
        .O(\memory_controller_inst/memory_controller_out_b [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[31]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [31]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[31]),
        .O(\memory_controller_inst/memory_controller_out_b [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[3]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [3]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[3]),
        .O(\memory_controller_inst/memory_controller_out_b [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[4]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [4]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[4]),
        .O(\memory_controller_inst/memory_controller_out_b [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[5]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [5]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[5]),
        .O(\memory_controller_inst/memory_controller_out_b [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[6]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [6]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[6]),
        .O(\memory_controller_inst/memory_controller_out_b [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[7]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [7]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[7]),
        .O(\memory_controller_inst/memory_controller_out_b [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[8]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [8]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[8]),
        .O(\memory_controller_inst/memory_controller_out_b [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h8F88)) 
    \memory_controller_out_reg_b[9]_i_1 
       (.I0(\memory_controller_inst/float_exception_flags/q_b_wire [9]),
        .I1(\memory_controller_inst/select_float_exception_flags_reg_b ),
        .I2(\memory_controller_inst/memory_controller_enable_reg_b ),
        .I3(memory_controller_out_b[9]),
        .O(\memory_controller_inst/memory_controller_out_b [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_1
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_34_n_0),
        .O(ram_reg_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_10
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_43_n_0),
        .O(ram_reg_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_11
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_44_n_0),
        .O(ram_reg_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_12
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_45_n_0),
        .O(ram_reg_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_13
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_46_n_0),
        .O(ram_reg_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_14
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_47_n_0),
        .O(ram_reg_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_15
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_48_n_0),
        .O(ram_reg_i_15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_16
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_49_n_0),
        .O(ram_reg_i_16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_17
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_50_n_0),
        .O(ram_reg_i_17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_18
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_51_n_0),
        .O(ram_reg_i_18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_19
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_52_n_0),
        .O(ram_reg_i_19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_2
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_35_n_0),
        .O(ram_reg_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_20
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_53_n_0),
        .O(ram_reg_i_20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_21
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_54_n_0),
        .O(ram_reg_i_21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_22
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_55_n_0),
        .O(ram_reg_i_22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_23
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_56_n_0),
        .O(ram_reg_i_23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_24
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_57_n_0),
        .O(ram_reg_i_24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_25
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_58_n_0),
        .O(ram_reg_i_25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_26
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_59_n_0),
        .O(ram_reg_i_26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_27
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_60_n_0),
        .O(ram_reg_i_27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000800082800000)) 
    ram_reg_i_28
       (.I0(ram_reg_i_61_n_0),
        .I1(\main_inst/cur_state_reg ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_memory_controller_in_a [4]),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .O(memory_controller_in_a));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_29
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_63_n_0),
        .O(ram_reg_i_29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_3
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_36_n_0),
        .O(ram_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_30
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_64_n_0),
        .O(ram_reg_i_30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_31
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_65_n_0),
        .O(ram_reg_i_31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_32
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_66_n_0),
        .O(ram_reg_i_32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00080000)) 
    ram_reg_i_33
       (.I0(ram_reg_i_67_n_0),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\select_float_exception_flags_reg_a[1]_i_1_n_0 ),
        .O(\memory_controller_inst/float_exception_flags_write_enable_a ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_34
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [31]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[31]),
        .O(ram_reg_i_34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_35
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [30]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[30]),
        .O(ram_reg_i_35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_36
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [29]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[29]),
        .O(ram_reg_i_36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_37
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [28]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[28]),
        .O(ram_reg_i_37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_38
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [27]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[27]),
        .O(ram_reg_i_38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_39
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [26]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[26]),
        .O(ram_reg_i_39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_4
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_37_n_0),
        .O(ram_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_40
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [25]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[25]),
        .O(ram_reg_i_40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_41
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [24]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[24]),
        .O(ram_reg_i_41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_42
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [23]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[23]),
        .O(ram_reg_i_42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_43
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [22]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[22]),
        .O(ram_reg_i_43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_44
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [21]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[21]),
        .O(ram_reg_i_44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_45
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [20]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[20]),
        .O(ram_reg_i_45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_46
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [19]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[19]),
        .O(ram_reg_i_46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_47
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [18]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[18]),
        .O(ram_reg_i_47_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_48
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [17]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[17]),
        .O(ram_reg_i_48_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_49
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [16]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[16]),
        .O(ram_reg_i_49_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_5
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_38_n_0),
        .O(ram_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_50
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [15]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[15]),
        .O(ram_reg_i_50_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_51
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [14]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[14]),
        .O(ram_reg_i_51_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_52
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [13]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[13]),
        .O(ram_reg_i_52_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_53
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [12]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[12]),
        .O(ram_reg_i_53_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_54
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [11]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[11]),
        .O(ram_reg_i_54_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_55
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [10]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[10]),
        .O(ram_reg_i_55_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_56
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [9]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[9]),
        .O(ram_reg_i_56_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_57
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [8]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[8]),
        .O(ram_reg_i_57_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_58
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [7]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[7]),
        .O(ram_reg_i_58_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_59
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [6]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[6]),
        .O(ram_reg_i_59_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_6
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_39_n_0),
        .O(ram_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_60
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [5]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[5]),
        .O(ram_reg_i_60_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    ram_reg_i_61
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[4] ),
        .O(ram_reg_i_61_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_62
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[4]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_63
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [3]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[3]),
        .O(ram_reg_i_63_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_64
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [2]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[2]),
        .O(ram_reg_i_64_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_65
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [1]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[1]),
        .O(ram_reg_i_65_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h9BFFFFBFDFFFFFBF)) 
    ram_reg_i_66
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_in_a [0]),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(memory_controller_out_a[0]),
        .O(ram_reg_i_66_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h64000040)) 
    ram_reg_i_67
       (.I0(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_write_enable_a ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg ),
        .O(ram_reg_i_67_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_68
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[31]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_69
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[30]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_7
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_40_n_0),
        .O(ram_reg_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_70
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[29]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_71
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[28]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_72
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[27]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_73
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[26]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_74
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[25]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_75
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[24]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_76
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[23]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_77
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[22]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_78
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[21]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_79
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[20]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_8
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_41_n_0),
        .O(ram_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_80
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[19]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_81
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[18]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_82
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[17]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_83
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[16]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_84
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[15]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_85
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[14]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_86
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[13]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_87
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[12]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_88
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[11]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_89
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[10]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0010)) 
    ram_reg_i_9
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(ram_reg_i_42_n_0),
        .O(ram_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_90
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[9]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_91
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[8]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_92
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[7]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_93
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[6]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_94
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[5]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000005004040)) 
    ram_reg_i_95
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(memory_controller_out_a[3]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040004)) 
    ram_reg_i_96
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[2]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000014040000)) 
    ram_reg_i_97
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(memory_controller_out_a[1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000005005040)) 
    ram_reg_i_98
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(memory_controller_out_a[0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_in_a [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00001044)) 
    ram_reg_i_99
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64_memory_controller_write_enable_a ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    \return_val[31]_i_1 
       (.I0(\return_val[31]_i_3_n_0 ),
        .I1(\return_val[31]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\return_val[31]_i_5_n_0 ),
        .O(\return_val[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0001000000000000)) 
    \return_val[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\return_val[31]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\return_val[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \return_val[31]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\return_val[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \return_val[31]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .O(\return_val[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF7FFFFFFFFFFFF)) 
    \return_val[31]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\return_val[31]_i_7_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\return_val[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \return_val[31]_i_6 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .O(\return_val[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \return_val[31]_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_[5] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\return_val[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000001)) 
    \return_val[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\return_val[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00010000)) 
    \return_val[63]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\return_val[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000002)) 
    \roundAndPackFloat64_0_1_reg[9]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFEF00000020)) 
    \roundAndPackFloat64_11_16_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSign_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\roundAndPackFloat64_11_16_reg[63]_i_2_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_11_16_reg ),
        .O(roundAndPackFloat64_11_16_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \roundAndPackFloat64_11_16_reg[63]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .O(\roundAndPackFloat64_11_16_reg[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFA6)) 
    \roundAndPackFloat64_57_0_reg[52]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [52]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [52]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_57_0_reg ),
        .O(roundAndPackFloat64_57_0_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8AAAAAAAAAAAAAA)) 
    \roundAndPackFloat64_57_0_reg[55]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [53]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hA8AAAAAAAAAAAAAA)) 
    \roundAndPackFloat64_57_0_reg[55]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [52]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[55]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [55]),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[55]_i_5 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [54]),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFA6)) 
    \roundAndPackFloat64_57_0_reg[55]_i_6 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [53]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [53]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_57_0_reg ),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFA6)) 
    \roundAndPackFloat64_57_0_reg[55]_i_7 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [52]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [52]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_57_0_reg ),
        .O(\roundAndPackFloat64_57_0_reg[55]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[59]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [59]),
        .O(\roundAndPackFloat64_57_0_reg[59]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[59]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [58]),
        .O(\roundAndPackFloat64_57_0_reg[59]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[59]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [57]),
        .O(\roundAndPackFloat64_57_0_reg[59]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[59]_i_5 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [56]),
        .O(\roundAndPackFloat64_57_0_reg[59]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10080000)) 
    \roundAndPackFloat64_57_0_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF9A009A)) 
    \roundAndPackFloat64_57_0_reg[63]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55_reg [63]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [63]),
        .I3(\main_inst/roundAndPackFloat64_57_0_reg ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_11_16_reg ),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[63]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [62]),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[63]_i_5 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [61]),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1000FFFF10001000)) 
    \roundAndPackFloat64_57_0_reg[63]_i_6 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg_reg_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_op_reg [60]),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h8)) 
    \roundAndPackFloat64_57_0_reg[63]_i_7 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .O(\roundAndPackFloat64_57_0_reg[63]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_57_0_reg_reg[55]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO(roundAndPackFloat64_57_0_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\roundAndPackFloat64_57_0_reg[55]_i_2_n_0 ,\roundAndPackFloat64_57_0_reg[55]_i_3_n_0 }),
        .O({\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_4 ,\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_5 ,\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_6 ,\roundAndPackFloat64_57_0_reg_reg[55]_i_1_n_7 }),
        .S({\roundAndPackFloat64_57_0_reg[55]_i_4_n_0 ,\roundAndPackFloat64_57_0_reg[55]_i_5_n_0 ,\roundAndPackFloat64_57_0_reg[55]_i_6_n_0 ,\roundAndPackFloat64_57_0_reg[55]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_57_0_reg_reg[59]_i_1 
       (.CI(roundAndPackFloat64_57_0_reg_reg[3]),
        .CO({\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_0 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_1 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_2 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_4 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_5 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_6 ,\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_7 }),
        .S({\roundAndPackFloat64_57_0_reg[59]_i_2_n_0 ,\roundAndPackFloat64_57_0_reg[59]_i_3_n_0 ,\roundAndPackFloat64_57_0_reg[59]_i_4_n_0 ,\roundAndPackFloat64_57_0_reg[59]_i_5_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_57_0_reg_reg[63]_i_2 
       (.CI(\roundAndPackFloat64_57_0_reg_reg[59]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_4 ,\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_5 ,\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_6 ,\roundAndPackFloat64_57_0_reg_reg[63]_i_2_n_7 }),
        .S({\roundAndPackFloat64_57_0_reg[63]_i_3_n_0 ,\roundAndPackFloat64_57_0_reg[63]_i_4_n_0 ,\roundAndPackFloat64_57_0_reg[63]_i_5_n_0 ,\roundAndPackFloat64_57_0_reg[63]_i_6_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(roundAndPackFloat64_arg_zExp),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [0]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[0]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [0]),
        .O(roundAndPackFloat64_arg_zExp));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[10]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[10]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [10]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[10]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [10]),
        .O(\roundAndPackFloat64_arg_zExp[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[11]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[11]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [11]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[11]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [11]),
        .O(\roundAndPackFloat64_arg_zExp[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[11]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[11]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[10] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[11]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[11]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[9] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[11]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[11]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[8] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[11]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[12]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[12]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [12]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[12]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [12]),
        .O(\roundAndPackFloat64_arg_zExp[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[13]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[13]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [13]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[13]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [13]),
        .O(\roundAndPackFloat64_arg_zExp[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[14]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[14]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [14]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[14]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [14]),
        .O(\roundAndPackFloat64_arg_zExp[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[15]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[15]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [15]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[15]_i_10 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[11]),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[15]_i_11 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[10]),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[15]_i_12 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[9]),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[15]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [15]),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[15]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[15]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[15]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[15]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[15]_i_9 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[12]),
        .O(\roundAndPackFloat64_arg_zExp[15]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[16]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[16]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [16]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[16]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [16]),
        .O(\roundAndPackFloat64_arg_zExp[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[17]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[17]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [17]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[17]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [17]),
        .O(\roundAndPackFloat64_arg_zExp[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[18]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[18]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [18]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[18]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [18]),
        .O(\roundAndPackFloat64_arg_zExp[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[19]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[19]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [19]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[19]_i_10 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[15]),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[19]_i_11 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[14]),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[19]_i_12 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[13]),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[19]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [19]),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[19]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[19]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[19]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[19]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[19]_i_9 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[16]),
        .O(\roundAndPackFloat64_arg_zExp[19]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[1]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[1]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [1]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[1]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [1]),
        .O(\roundAndPackFloat64_arg_zExp[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[20]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[20]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [20]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[20]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [20]),
        .O(\roundAndPackFloat64_arg_zExp[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[21]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[21]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [21]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[21]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [21]),
        .O(\roundAndPackFloat64_arg_zExp[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[22]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[22]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [22]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[22]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [22]),
        .O(\roundAndPackFloat64_arg_zExp[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[23]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[23]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [23]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[23]_i_10 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[19]),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[23]_i_11 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[18]),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[23]_i_12 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[17]),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[23]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [23]),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[23]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[23]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[23]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[23]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[23]_i_9 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[20]),
        .O(\roundAndPackFloat64_arg_zExp[23]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[24]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[24]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [24]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[24]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [24]),
        .O(\roundAndPackFloat64_arg_zExp[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[25]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[25]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [25]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[25]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [25]),
        .O(\roundAndPackFloat64_arg_zExp[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[26]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[26]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [26]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[26]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [26]),
        .O(\roundAndPackFloat64_arg_zExp[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[27]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[27]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [27]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[27]_i_10 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[23]),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[27]_i_11 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[22]),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[27]_i_12 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[21]),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[27]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [27]),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[27]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[27]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[27]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[27]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[27]_i_9 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[24]),
        .O(\roundAndPackFloat64_arg_zExp[27]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[28]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[28]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [28]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[28]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [28]),
        .O(\roundAndPackFloat64_arg_zExp[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[29]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[29]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [29]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[29]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [29]),
        .O(\roundAndPackFloat64_arg_zExp[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[2]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[2]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [2]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[2]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [2]),
        .O(\roundAndPackFloat64_arg_zExp[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[30]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[30]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [30]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[30]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [30]),
        .O(\roundAndPackFloat64_arg_zExp[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[31]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [31]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_10 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[31]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_11 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[30]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_12 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[29]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_13 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[28]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_14 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[27]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_15 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[26]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[31]_i_16 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[25]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[31]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [31]),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[31]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[31]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[31]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[31]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[31]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[3]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[3]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [3]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[3]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [3]),
        .O(\roundAndPackFloat64_arg_zExp[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[3]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[3]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[2] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[3]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[3]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zExp[3]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[0]),
        .O(\roundAndPackFloat64_arg_zExp[3]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[4]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[4]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [4]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[4]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [4]),
        .O(\roundAndPackFloat64_arg_zExp[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[5]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[5]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [5]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[5]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [5]),
        .O(\roundAndPackFloat64_arg_zExp[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[6]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[6]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [6]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[6]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_5 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [6]),
        .O(\roundAndPackFloat64_arg_zExp[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[7]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[7]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [7]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[7]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_4 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [7]),
        .O(\roundAndPackFloat64_arg_zExp[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[7]_i_4 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[7] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_5 ),
        .O(\roundAndPackFloat64_arg_zExp[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[7]_i_5 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[6] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_6 ),
        .O(\roundAndPackFloat64_arg_zExp[7]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[7]_i_6 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[5] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zExp[7]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \roundAndPackFloat64_arg_zExp[7]_i_7 
       (.I0(\main_inst/main_195_196_reg_reg_n_0_[4] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zExp[7]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[8]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[8]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [8]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[8]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_7 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [8]),
        .O(\roundAndPackFloat64_arg_zExp[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zExp[9]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zExp[9]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zExp1ii_reg [9]),
        .O(\main_inst/roundAndPackFloat64_arg_zExp [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEF0040)) 
    \roundAndPackFloat64_arg_zExp[9]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_6 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/main_101_zExp1ii_reg [9]),
        .O(\roundAndPackFloat64_arg_zExp[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[11]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_0 ),
        .CO(roundAndPackFloat64_arg_zExp_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[10] ,\main_inst/main_195_196_reg_reg_n_0_[9] ,\main_inst/main_195_196_reg_reg_n_0_[8] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[11]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[11]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[11]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[11]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[11]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[15]_i_3 
       (.CI(roundAndPackFloat64_arg_zExp_reg[3]),
        .CO({\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[15]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[15]_i_8 
       (.CI(roundAndPackFloat64_arg_zSig_reg[3]),
        .CO({\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_0 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_1 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_2 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_4 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_5 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_6 ,\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[15]_i_9_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_10_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_11_n_0 ,\roundAndPackFloat64_arg_zExp[15]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[19]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[15]_i_3_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[19]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[19]_i_8 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[15]_i_8_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_0 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_1 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_2 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_4 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_5 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_6 ,\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[19]_i_9_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_10_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_11_n_0 ,\roundAndPackFloat64_arg_zExp[19]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[23]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[19]_i_3_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[23]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[23]_i_8 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[19]_i_8_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_0 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_1 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_2 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_4 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_5 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_6 ,\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[23]_i_9_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_10_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_11_n_0 ,\roundAndPackFloat64_arg_zExp[23]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[27]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[23]_i_3_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[27]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[27]_i_8 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[23]_i_8_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_0 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_1 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_2 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_4 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_5 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_6 ,\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[27]_i_9_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_10_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_11_n_0 ,\roundAndPackFloat64_arg_zExp[27]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[31]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[27]_i_3_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] ,\main_inst/main_195_196_reg_reg_n_0_[31] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[31]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[31]_i_8 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_4 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_5 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_6 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_8_n_7 }),
        .S({\<const0>__0__0 ,\roundAndPackFloat64_arg_zExp[31]_i_10_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_11_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[31]_i_9 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[27]_i_8_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_0 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_1 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_2 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_4 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_5 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_6 ,\roundAndPackFloat64_arg_zExp_reg[31]_i_9_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[31]_i_13_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_14_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_15_n_0 ,\roundAndPackFloat64_arg_zExp[31]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[3]_i_3 
       (.CI(\<const0>__0__0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_3 }),
        .CYINIT(\<const1>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[3] ,\main_inst/main_195_196_reg_reg_n_0_[2] ,\main_inst/main_195_196_reg_reg_n_0_[1] ,\main_inst/main_195_196_reg_reg_n_0_ }),
        .O({\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[3]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[3]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[3]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[3]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zExp_reg[7]_i_3 
       (.CI(\roundAndPackFloat64_arg_zExp_reg[3]_i_3_n_0 ),
        .CO({\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_0 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_1 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_2 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_195_196_reg_reg_n_0_[7] ,\main_inst/main_195_196_reg_reg_n_0_[6] ,\main_inst/main_195_196_reg_reg_n_0_[5] ,\main_inst/main_195_196_reg_reg_n_0_[4] }),
        .O({\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_4 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_5 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_6 ,\roundAndPackFloat64_arg_zExp_reg[7]_i_3_n_7 }),
        .S({\roundAndPackFloat64_arg_zExp[7]_i_4_n_0 ,\roundAndPackFloat64_arg_zExp[7]_i_5_n_0 ,\roundAndPackFloat64_arg_zExp[7]_i_6_n_0 ,\roundAndPackFloat64_arg_zExp[7]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[0]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(roundAndPackFloat64_arg_zSig),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    \roundAndPackFloat64_arg_zSig[0]_i_2 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zSig[1]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .O(roundAndPackFloat64_arg_zSig));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[10]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[10]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_ ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[10]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[11]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[10]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_ ),
        .O(\roundAndPackFloat64_arg_zSig[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[10]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[10]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[12]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \roundAndPackFloat64_arg_zSig[10]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .O(\roundAndPackFloat64_arg_zSig[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[11]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[11]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[11] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[11]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[12]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[11]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[11] ),
        .O(\roundAndPackFloat64_arg_zSig[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[11]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[11]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[13]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \roundAndPackFloat64_arg_zSig[11]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[15]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[12]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[12]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[12] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[12]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[13]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[12]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[12] ),
        .O(\roundAndPackFloat64_arg_zSig[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[12]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[12]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[14]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \roundAndPackFloat64_arg_zSig[12]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[16]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[13]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[13]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[13] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[13]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[14]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[13]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[13] ),
        .O(\roundAndPackFloat64_arg_zSig[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_arg_zSig[13]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[15]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[13]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \roundAndPackFloat64_arg_zSig[13]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[17]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[14]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[14]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[14] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[14]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[15]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[14]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[14] ),
        .O(\roundAndPackFloat64_arg_zSig[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_arg_zSig[14]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[16]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[14]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0004FFFF00040000)) 
    \roundAndPackFloat64_arg_zSig[14]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[18]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[15]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[15]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[15] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[15]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[16]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[15]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[15] ),
        .O(\roundAndPackFloat64_arg_zSig[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[15]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[15]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[17]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[15]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[16]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[16]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[16] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[16]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[17]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[16]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[16] ),
        .O(\roundAndPackFloat64_arg_zSig[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[16]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[16]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[18]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[16]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[17]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[17]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[17] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[17]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[18]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[17]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[17] ),
        .O(\roundAndPackFloat64_arg_zSig[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[17]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[17]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[17]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[18]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[18]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[18] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[18]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[19]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[18]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[18] ),
        .O(\roundAndPackFloat64_arg_zSig[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[18]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[18]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[18]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[19]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[19]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[19] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[19]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[20]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[19]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[19] ),
        .O(\roundAndPackFloat64_arg_zSig[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[19]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[19]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[1]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[1]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[1] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[1]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[2]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[1]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_arg_zSig[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \roundAndPackFloat64_arg_zSig[1]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[20]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[20]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[20] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[20]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[21]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[20]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[20] ),
        .O(\roundAndPackFloat64_arg_zSig[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[20]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[20]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[20]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[21]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[21]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[21] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[21]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[22]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[21]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[21] ),
        .O(\roundAndPackFloat64_arg_zSig[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[21]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[21]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[21]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[22]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[22]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[22] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[22]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[23]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[22]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[22] ),
        .O(\roundAndPackFloat64_arg_zSig[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[22]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000B08)) 
    \roundAndPackFloat64_arg_zSig[22]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .O(\roundAndPackFloat64_arg_zSig[22]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[23]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[23]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[23] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[23]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[24]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[23]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[23] ),
        .O(\roundAndPackFloat64_arg_zSig[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[23]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[23]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[23]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[24]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[24]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[24] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[24]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[25]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[24]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[24] ),
        .O(\roundAndPackFloat64_arg_zSig[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[24]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I3(\roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I5(\roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[24]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[25]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[25]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[25] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[25]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[26]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[25]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[25] ),
        .O(\roundAndPackFloat64_arg_zSig[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[25]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[25]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[26]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[26]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[26] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[26]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[27]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[26]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[26] ),
        .O(\roundAndPackFloat64_arg_zSig[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[26]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[26]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[27]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[27]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[27] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[27]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[28]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[27]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[27] ),
        .O(\roundAndPackFloat64_arg_zSig[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[27]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[27]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[28]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[28]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[28] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[28]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[29]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[28]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[28] ),
        .O(\roundAndPackFloat64_arg_zSig[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[28]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[28]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[29]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[29]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[29] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[29]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[30]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[29]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[29] ),
        .O(\roundAndPackFloat64_arg_zSig[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[29]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[29]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[2]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[2]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[2] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[2]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[3]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[2]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000010)) 
    \roundAndPackFloat64_arg_zSig[2]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[2]_i_5 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[8]),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[2]_i_6 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[7]),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[2]_i_7 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ),
        .I1(memory_controller_out_a[6]),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[2]_i_8 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[5] ),
        .I1(memory_controller_out_a[5]),
        .O(\roundAndPackFloat64_arg_zSig[2]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[30]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[30]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[30] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[30]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[31]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[30]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[30] ),
        .O(\roundAndPackFloat64_arg_zSig[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[30]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000030BB3088)) 
    \roundAndPackFloat64_arg_zSig[30]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[31]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[31]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[31] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[31]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[32]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[31]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[31] ),
        .O(\roundAndPackFloat64_arg_zSig[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[31]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[31]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[31]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[31]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[31]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[32]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[32]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[32] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[32]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[33]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[32]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[32] ),
        .O(\roundAndPackFloat64_arg_zSig[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[32]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[32]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[32]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[32]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[32]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[33]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[33]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[33] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[33]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[34]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[33]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[33] ),
        .O(\roundAndPackFloat64_arg_zSig[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[33]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[33]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[33]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[33]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[33]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[33]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[34]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[34]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[34] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[34]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[35]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[34]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[34] ),
        .O(\roundAndPackFloat64_arg_zSig[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[34]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[34]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[34]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[34]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[34]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[34]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[35]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[35]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[35] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[35]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[36]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[35]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[35] ),
        .O(\roundAndPackFloat64_arg_zSig[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[35]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[35]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[35]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[35]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[35]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[35]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[36]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[36]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[36] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[36]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[37]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[36]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[36] ),
        .O(\roundAndPackFloat64_arg_zSig[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[36]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[36]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[36]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[36]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[36]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[36]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[37]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[37]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[37] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[37]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[38]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[37]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[37] ),
        .O(\roundAndPackFloat64_arg_zSig[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[37]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[37]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[37]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[37]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[37]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[38]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[38]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[38] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[38]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[39]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[38]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[38] ),
        .O(\roundAndPackFloat64_arg_zSig[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[38]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[38]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[38]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00B8)) 
    \roundAndPackFloat64_arg_zSig[38]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[38]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[39]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[39]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[39] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[39]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[40]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[39]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[39] ),
        .O(\roundAndPackFloat64_arg_zSig[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[39]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[39]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[47]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[3]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[3]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[3] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[3]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[4]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[3]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_arg_zSig[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[3]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[3]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[5]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \roundAndPackFloat64_arg_zSig[3]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .O(\roundAndPackFloat64_arg_zSig[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[40]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[40]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[40] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[40]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[41]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[40]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[40] ),
        .O(\roundAndPackFloat64_arg_zSig[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[40]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[40]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[40]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[48]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[40]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[41]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[41]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[41] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[41]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[42]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[41]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_arg_zSig[41]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[41]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[43]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[41]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[49]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[41]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[42]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[42]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[42] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[42]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[43]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[42]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[42] ),
        .O(\roundAndPackFloat64_arg_zSig[42]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_arg_zSig[42]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[44]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[42]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[42]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[50]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[42]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[43]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[43]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[43] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[43]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[44]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[43]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[43] ),
        .O(\roundAndPackFloat64_arg_zSig[43]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[43]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[45]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[43]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[43]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[43]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[51]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[43]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[43]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[47]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[43]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[44]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[44]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[44] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[44]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[45]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[44]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[44] ),
        .O(\roundAndPackFloat64_arg_zSig[44]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[44]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[46]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[44]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[44]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[44]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[52]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[44]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[44]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[48]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[44]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[45]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[45]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[45]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[46]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[45]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[45]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_arg_zSig[45]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[45]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig[47]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[45]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[45]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[53]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[45]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[45]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[49]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[45]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[46]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[46]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[46]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[47]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[46]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[46]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_arg_zSig[46]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[46]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig[48]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[46]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00B8FFFF00B80000)) 
    \roundAndPackFloat64_arg_zSig[46]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[54]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[46]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[46]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[50]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[46]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[47]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[47]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[47]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[48]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[47]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[47]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[47]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[47]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[49]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[47]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[47]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[47]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[51]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[47]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[47]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ),
        .O(\roundAndPackFloat64_arg_zSig[47]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[48]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[48]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[48]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[49]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[48]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[48]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[48]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[48]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[50]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[48]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[48]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[48]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[52]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[48]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[48]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ),
        .O(\roundAndPackFloat64_arg_zSig[48]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[49]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[49]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[49]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[50]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[49]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[49]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[49]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[51]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[49]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[49]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[49]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[53]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[49]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[49]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[34] ),
        .O(\roundAndPackFloat64_arg_zSig[49]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[4]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[4]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[4] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[4]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[5]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[4]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_arg_zSig[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[4]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[4]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[6]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \roundAndPackFloat64_arg_zSig[4]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .O(\roundAndPackFloat64_arg_zSig[4]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[50]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[50]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[50]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[51]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[50]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[50]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[50]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[50]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[52]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[50]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[50]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[50]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[54]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[50]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[50]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[35] ),
        .O(\roundAndPackFloat64_arg_zSig[50]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[51]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[51]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[51]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[52]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[51]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[51]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[51]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[51]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[53]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[51]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[51]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[51]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[59]_i_7_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[51]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[51]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[36] ),
        .O(\roundAndPackFloat64_arg_zSig[51]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[52]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[52]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[52]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[53]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[52]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[52]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[52]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[52]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[54]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[52]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[52]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[52]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[60]_i_7_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[52]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[52]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[37] ),
        .O(\roundAndPackFloat64_arg_zSig[52]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[53]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[53]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[53]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[54]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[53]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[53]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[53]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[55]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[53]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[53]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[53]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[61]_i_7_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[53]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[53]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[38] ),
        .O(\roundAndPackFloat64_arg_zSig[53]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[54]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[54]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[54]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[55]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[54]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[54]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[54]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[54]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[56]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[54]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[54]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[54]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[54]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[54]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[39] ),
        .O(\roundAndPackFloat64_arg_zSig[54]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[55]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[55]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[55]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[56]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[55]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[55]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[55]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[55]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[57]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[55]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[55]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[59]_i_7_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[63]_i_19_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[55]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[55]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ),
        .O(\roundAndPackFloat64_arg_zSig[55]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[56]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[56]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[56]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[57]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[56]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[56]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[56]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[56]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[58]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[56]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[56]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[60]_i_7_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[63]_i_11_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[56]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[56]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_arg_zSig[56]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[57]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[57]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[57]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[58]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[57]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_arg_zSig[57]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[59]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[59]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[57]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[57]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[61]_i_7_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[63]_i_21_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[57]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[57]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ),
        .O(\roundAndPackFloat64_arg_zSig[57]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[58]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[58]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[58]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[59]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[58]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[58]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_arg_zSig[58]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[60]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[60]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[58]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[58]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[58]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[62]_i_7_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I3(\roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I5(\roundAndPackFloat64_arg_zSig[63]_i_17_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[58]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[58]_i_5 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ),
        .O(\roundAndPackFloat64_arg_zSig[58]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[59]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[59]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[59]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[60]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[59]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[59]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[61]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[61]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[59]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[59]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[59]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_19_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[59]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[59]_i_7_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[59]_i_8_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[59]_i_6 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[59]_i_7 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[32] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[16] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[48] ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[59]_i_8 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[8] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[40] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[24] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[56] ),
        .O(\roundAndPackFloat64_arg_zSig[59]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[5]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[5]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[5] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[5]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[6]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[5]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_arg_zSig[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[5]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[5]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[7]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \roundAndPackFloat64_arg_zSig[5]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .O(\roundAndPackFloat64_arg_zSig[5]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[60]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[60]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[60]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[61]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[60]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF33CC00B8B8B8B8)) 
    \roundAndPackFloat64_arg_zSig[60]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[62]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[62]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig[60]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_arg_zSig[60]_i_5_n_0 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[60]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_11_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[60]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[60]_i_7_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[60]_i_8_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[60]_i_6 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[60]_i_7 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[33] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[17] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[49] ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[60]_i_8 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[9] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[41] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[25] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[57] ),
        .O(\roundAndPackFloat64_arg_zSig[60]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10000000)) 
    \roundAndPackFloat64_arg_zSig[61]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[61]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h45400000)) 
    \roundAndPackFloat64_arg_zSig[61]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[62]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[61]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_arg_zSig[61]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[61]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[61]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_9_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[61]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_21_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[61]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[61]_i_7_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[61]_i_8_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[61]_i_6 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[61]_i_7 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[34] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[18] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[50] ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[61]_i_8 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[10] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[42] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[26] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[58] ),
        .O(\roundAndPackFloat64_arg_zSig[61]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[62]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[62]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[62] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[62]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[63]_i_5_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[62]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[62] ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_arg_zSig[62]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[62]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[62]_i_5_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_6_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[62]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_17_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[62]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[62]_i_7_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I2(\roundAndPackFloat64_arg_zSig[62]_i_8_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_arg_zSig[62]_i_6 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I4(\main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[62]_i_7 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[35] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[19] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[51] ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[62]_i_8 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[11] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[43] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[27] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[59] ),
        .O(\roundAndPackFloat64_arg_zSig[62]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[63]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[63] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_arg_zSig[63]_i_10 
       (.I0(\roundAndPackFloat64_arg_zSig[61]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_21_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_22_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_11 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[37] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[21] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[53] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_12 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[13] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[45] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[29] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[61] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[63]_i_13 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[4] ),
        .I1(memory_controller_out_a[4]),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h6)) 
    \roundAndPackFloat64_arg_zSig[63]_i_14 
       (.I0(\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[3] ),
        .I1(memory_controller_out_a[3]),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \roundAndPackFloat64_arg_zSig[63]_i_15 
       (.I0(memory_controller_out_a[2]),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \roundAndPackFloat64_arg_zSig[63]_i_16 
       (.I0(memory_controller_out_a[1]),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_17 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[7] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[39] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[23] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[55] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_18 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[15] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[47] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[31] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[63] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_19 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[36] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[20] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[52] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[63]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[63]_i_4_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[63]_i_5_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[63] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_20 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[12] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[44] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[28] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[60] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_21 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[38] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[22] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[54] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_arg_zSig[63]_i_22 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[14] ),
        .I1(\main_inst/main_195_zSig0ii_reg_reg_n_0_[46] ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[30] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\main_inst/main_195_zSig0ii_reg_reg_n_0_[62] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hEA)) 
    \roundAndPackFloat64_arg_zSig[63]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[63]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_6_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_8_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[63]_i_5 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_10_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_arg_zSig[63]_i_6 
       (.I0(\roundAndPackFloat64_arg_zSig[60]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_11_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_12_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_arg_zSig[63]_i_8 
       (.I0(\roundAndPackFloat64_arg_zSig[62]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_17_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_18_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_arg_zSig[63]_i_9 
       (.I0(\roundAndPackFloat64_arg_zSig[59]_i_5_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig[63]_i_19_n_0 ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I4(\roundAndPackFloat64_arg_zSig[63]_i_20_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[63]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[6]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[6]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[6]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[7]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[6]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[6] ),
        .O(\roundAndPackFloat64_arg_zSig[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[6]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[6]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[8]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000010)) 
    \roundAndPackFloat64_arg_zSig[6]_i_4 
       (.I0(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I2(\main_inst/main_195_zSig0ii_reg_reg_n_0_[3] ),
        .I3(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .O(\roundAndPackFloat64_arg_zSig[6]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[7]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[7]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[7] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[7]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[8]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[7]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[7] ),
        .O(\roundAndPackFloat64_arg_zSig[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[7]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[7]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[9]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \roundAndPackFloat64_arg_zSig[7]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_ ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[4] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .O(\roundAndPackFloat64_arg_zSig[7]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[8]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[8]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[8] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[8]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[9]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[8]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[8] ),
        .O(\roundAndPackFloat64_arg_zSig[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[8]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[8]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[10]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \roundAndPackFloat64_arg_zSig[8]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[5] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .O(\roundAndPackFloat64_arg_zSig[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFEFFFFFF10000000)) 
    \roundAndPackFloat64_arg_zSig[9]_i_1 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .I2(\roundAndPackFloat64_arg_zSig[9]_i_2_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[9] ),
        .O(\main_inst/roundAndPackFloat64_arg_zSig [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEFEAFFFF45400000)) 
    \roundAndPackFloat64_arg_zSig[9]_i_2 
       (.I0(\roundAndPackFloat64_arg_zSig[63]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig[10]_i_3_n_0 ),
        .I2(memory_controller_out_a[0]),
        .I3(\roundAndPackFloat64_arg_zSig[9]_i_3_n_0 ),
        .I4(main_1_4_reg),
        .I5(\main_inst/main_101_zSig0i12i_reg_reg_n_0_[9] ),
        .O(\roundAndPackFloat64_arg_zSig[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_arg_zSig[9]_i_3 
       (.I0(\roundAndPackFloat64_arg_zSig[9]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 ),
        .I2(\roundAndPackFloat64_arg_zSig[11]_i_4_n_0 ),
        .O(\roundAndPackFloat64_arg_zSig[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000B08)) 
    \roundAndPackFloat64_arg_zSig[9]_i_4 
       (.I0(\main_inst/main_195_zSig0ii_reg_reg_n_0_[2] ),
        .I1(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ),
        .I2(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ),
        .I3(\main_inst/main_195_zSig0ii_reg_reg_n_0_[6] ),
        .I4(\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 ),
        .I5(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ),
        .O(\roundAndPackFloat64_arg_zSig[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zSig_reg[2]_i_4 
       (.CI(\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_0 ),
        .CO(roundAndPackFloat64_arg_zSig_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_ ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[5] }),
        .O({\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_4 ,\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_5 ,\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_6 ,\roundAndPackFloat64_arg_zSig_reg[2]_i_4_n_7 }),
        .S({\roundAndPackFloat64_arg_zSig[2]_i_5_n_0 ,\roundAndPackFloat64_arg_zSig[2]_i_6_n_0 ,\roundAndPackFloat64_arg_zSig[2]_i_7_n_0 ,\roundAndPackFloat64_arg_zSig[2]_i_8_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_arg_zSig_reg[63]_i_7 
       (.CI(\<const0>__0__0 ),
        .CO({\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_0 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_1 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_2 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_3 }),
        .CYINIT(memory_controller_out_a[0]),
        .DI({\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[4] ,\main_inst/main_normalizeRoundAndPackFloat64exitii_209_reg_reg_n_0_[3] ,\<const1>__0__0 ,\<const1>__0__0 }),
        .O({\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_4 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_5 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_6 ,\roundAndPackFloat64_arg_zSig_reg[63]_i_7_n_7 }),
        .S({\roundAndPackFloat64_arg_zSig[63]_i_13_n_0 ,\roundAndPackFloat64_arg_zSig[63]_i_14_n_0 ,\roundAndPackFloat64_arg_zSig[63]_i_15_n_0 ,\roundAndPackFloat64_arg_zSig[63]_i_16_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hBAAAAAAAAAAAAAAA)) 
    \roundAndPackFloat64_arg_zSign[0]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_start ),
        .I1(\roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[6] ),
        .I4(\main_inst/cur_state_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_arg_zSign[0]_i_5_n_0 ),
        .O(\main_inst/roundAndPackFloat64_arg_zSign ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h2000000000000000)) 
    \roundAndPackFloat64_arg_zSign[0]_i_2 
       (.I0(\main_inst/main_195_0ii_reg ),
        .I1(\roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ),
        .I2(\roundAndPackFloat64_arg_zSign[0]_i_5_n_0 ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\main_inst/cur_state_reg_n_0_[6] ),
        .O(roundAndPackFloat64_arg_zSign));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000001000)) 
    \roundAndPackFloat64_arg_zSign[0]_i_3 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_1_scevgep_reg[31]_i_3_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\main_inst/roundAndPackFloat64_start ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \roundAndPackFloat64_arg_zSign[0]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_arg_zSign[0]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \roundAndPackFloat64_arg_zSign[0]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[2] ),
        .I1(\main_inst/cur_state_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_arg_zSign[0]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF000000A2)) 
    roundAndPackFloat64_finish_reg_i_1
       (.I0(\main_inst/roundAndPackFloat64_finish_reg_reg_n_0 ),
        .I1(\roundAndPackFloat64_return_val_reg[63]_i_4_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(reset),
        .I4(\main_inst/roundAndPackFloat64_finish_reg1 ),
        .I5(\main_inst/roundAndPackFloat64_finish ),
        .O(roundAndPackFloat64_finish_reg_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h32333232)) 
    \roundAndPackFloat64_return_val_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_finish_reg1 ),
        .I1(\main_inst/roundAndPackFloat64_finish ),
        .I2(reset),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_return_val_reg[63]_i_4_n_0 ),
        .O(roundAndPackFloat64_return_val_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFEFFFEFE)) 
    \roundAndPackFloat64_return_val_reg[63]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_finish_reg1 ),
        .I1(\main_inst/roundAndPackFloat64_finish ),
        .I2(reset),
        .I3(\main_inst/cur_state_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_return_val_reg[63]_i_4_n_0 ),
        .O(\roundAndPackFloat64_return_val_reg[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAAAAAAAABAA)) 
    \roundAndPackFloat64_return_val_reg[63]_i_3 
       (.I0(reset),
        .I1(\roundAndPackFloat64_return_val_reg[63]_i_5_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_shift64RightJammingexitii_z0iii_reg[41]_i_6_n_0 ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .I5(\main_inst/cur_state_reg_n_0_ ),
        .O(\main_inst/roundAndPackFloat64_finish_reg1 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000100)) 
    \roundAndPackFloat64_return_val_reg[63]_i_4 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[4] ),
        .I2(\main_inst/cur_state_reg_n_0_[6] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg_n_0_[2] ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_return_val_reg[63]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \roundAndPackFloat64_return_val_reg[63]_i_5 
       (.I0(\main_inst/cur_state_reg_n_0_[1] ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_return_val_reg[63]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \roundAndPackFloat64_shift64RightJammingexit_34_reg[9]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFACAFFFFFACA0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_31_33 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_3_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_2_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_21_29 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [0]),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_100 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ),
        .O(roundAndPackFloat64_shift64RightJammingexit_z0i_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_101 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_101_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_102 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_102_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_103 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_103_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_107 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_107_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_108 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_108_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_109 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_109_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h8FFF8F558FAA8F00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_11 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_25_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_26_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_27_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_110 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_110_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3202)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_112 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_124_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_154_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_155_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_112_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h005C00FF005C0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_113 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_158_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_155_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_113_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF005C0000005C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_114 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_159_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_160_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_114_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00005C5C0000FF00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_115 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_160_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_163_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_115_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_116 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_164_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_165_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_116_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_117 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_140_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_165_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_166_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_117_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_168_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_169_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_137_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF008F008F)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_12 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_25_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_28_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_29_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_120 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_164_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_166_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_170_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_120_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_121 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_170_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_171_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_172_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_121_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_122 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_173_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_172_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_122_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_123 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_173_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_171_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_174_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_175_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_123_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h553355330F000FFF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_124 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_124_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_125 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_179_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_125_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_126 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_126_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_127 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_129_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_127_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_128 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_128_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_129 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_129_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_132 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_132_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_133 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_181_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_133_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_134 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_138_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_132_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_134_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_135 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_182_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_179_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_135_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_136 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_183_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_181_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_136_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_137 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_184_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_137_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_138 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_138_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_139 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_185_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_139_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_14 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_140 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_186_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_182_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_140_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_144_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_146 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_146_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_147 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_147_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_148 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_148_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_149 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_149_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_15 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF005C0000005C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_150 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_187_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_188_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_150_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3202)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_151 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_188_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_189_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_190_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_151_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF03AA020000AA02)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_152 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_190_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_191_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_192_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_193_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_194_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_152_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFCFFFCFFF00FF0D)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_153 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_195_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_196_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_197_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_198_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_153_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_154 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_199_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_174_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_200_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_201_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_154_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_155 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_202_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_201_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_155_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB080FFFFB0800000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_204_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_158 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_202_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_200_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_205_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_157_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_158_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_159 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_156_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_205_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_206_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_207_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_159_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_16 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_160 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_208_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_207_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_160_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30BB000030880000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44FFFFCF77FFFF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_163 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_208_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_206_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_209_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_162_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_163_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_164 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_210_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_186_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_164_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_165 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_211_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_183_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_165_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_166 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_168_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_139_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_166_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_168 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_212_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_168_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_169 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_213_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_169_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_17 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_170 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_214_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_211_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_170_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_171 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_169_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_171_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_172 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_215_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_210_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_172_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_173 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_216_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_214_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_173_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_174 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_217_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_215_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_174_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_175 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_167_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_175_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_179 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_179_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_18 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_181 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_181_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_182 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_145_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_182_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_183 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_180_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_183_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_184 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_184_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_185 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_185_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_186 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_218_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_186_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_187 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_161_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_209_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_219_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_220_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_187_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h5C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_188 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_221_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_220_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_188_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF0EEFFEE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_189 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_221_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_219_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_192_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_222_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_189_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFF7FFF7FFFF0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_190 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_222_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_190_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAAAAAABAAAAAAAA)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_191 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_191_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_192 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_192_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCCC0CCC4CCCCCCCC)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_193 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_193_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFF4F7F)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_194 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_194_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_195 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_195_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h10)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_196 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_196_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_197 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_197_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h02)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_198 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_198_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_199 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_176_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_177_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_199_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00470047000000FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_20 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_42_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_29_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB080FFFFB0800000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_200 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_178_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_200_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_201 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_223_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_216_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_201_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB080FFFFB0800000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_202 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_217_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_202_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_204 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_204_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB080FFFFB0800000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_205 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_223_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_205_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB080FFFFB0800000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_206 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_224_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_206_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h4F7F00004F7FFFFF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_207 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_225_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_207_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB800FFFFB8000000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_208 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_226_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_208_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h30BB000030880000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_209 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_209_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF00004747)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_21 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_43_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_44_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_210 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_227_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_210_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_211 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_228_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_211_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_212 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_212_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_213 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_213_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00E2FFFF00E20000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_214 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_229_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_214_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_215 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_215_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_216 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_216_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_217 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_217_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_218 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_218_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_219 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_219_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00470047000000FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_22 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_47_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_43_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCF44CF77FFFFFFFF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_220 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_203_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_220_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000000000000B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_221 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_221_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_222 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_222_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000033B800B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_223 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_223_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_224 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_224_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_225 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_225_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000B0008)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_226 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_226_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_227 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_227_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_228 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_228_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h00E2)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_229 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_229_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF00004747)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_23 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_48_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_49_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h474700CC474733FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_51_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_53_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFEAEAAAAFEAE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_25 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_54_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_56_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h474700CC474733FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_26 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_58_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_60_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h474700CC474733FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_27 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_62_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_64_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF77F077)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_28 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_24_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_26_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_65_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_66_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_29 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_67_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_66_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hCFC0AFAFCFC0A0A0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_2_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_3_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_8_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_9_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_31 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_32 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_33 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_34 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h1103)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_36 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_78_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_79_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_48_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00004747000000FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_37 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_78_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_82_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF00470047)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_38 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_83_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_84_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00470047000000FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_39 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_87_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_84_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_51_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_42 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_67_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_65_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_92_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_41_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_43 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_93_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_94_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_44 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_40_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_92_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_95_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_94_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_47 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_93_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_95_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_99_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_46_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_48 
       (.I0(roundAndPackFloat64_shift64RightJammingexit_z0i_reg),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_101_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_48_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_49 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_45_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_99_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_102_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_101_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_49_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_51 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_51_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_53 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_53_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_54 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_54_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_56 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_103_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_56_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_58 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_58_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_6 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_60 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_60_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_62 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_62_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_64 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_64_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_65 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_55_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_56_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_65_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_66 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_62_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_66_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hB8B8B8B8FF33CC00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_67 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_58_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_67_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_69 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_69_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_7 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_70 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_70_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_71 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_71_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h01)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_72 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_72_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000000FF00004747)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_74 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_116_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_117_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_74_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00005C5C000000FF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_75 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_116_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_120_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_75_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FF005C0000005C)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_76 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_118_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_119_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_121_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_122_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_76_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h3202)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_77 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_122_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_123_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_124_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_77_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_78 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_125_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_126_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_78_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_79 
       (.I0(roundAndPackFloat64_shift64RightJammingexit_z0i_reg),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_102_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_126_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_127_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_79_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_8 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_128_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_129_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFF00B8B8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_130_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_132_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_82 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_125_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_127_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_81_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_133_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_82_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_83 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_80_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_133_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_134_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_135_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_83_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_84 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_136_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_135_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_84_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_137_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_138_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_85_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_139_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_128_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFEEF0EE)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_87 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_136_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_134_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_140_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_86_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_87_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_88_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_89_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_9 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_3_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_18_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_90_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_92 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_63_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_92_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_93 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_142_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_104_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_141_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_61_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_93_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_94 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_59_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_94_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_95 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_50_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_91_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_52_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_95_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_96_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_97_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h30BB3088)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_98_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_99 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_143_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_105_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_131_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_57_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_99_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hD1FFD100)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22222228EEEEEEEB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8BFF8B00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7777777D44444441)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB888B8BB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB888B8BB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF5F503F3)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hBB8B888B)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB888B8BB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF5F503F3)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[18]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[19]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00D8FFD8)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_2_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_3_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8FFB800)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_3_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_5_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFAFCFC0A0A0CFC0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_5 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[20]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[21]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[22]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[23]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF5F503F3)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[24]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[25]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[26]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[27]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[28]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[29]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28E82BEB282BE8EB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_4_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_5_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_4 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_5 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[2]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[30]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[31]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFF47FFFFFF470000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[32]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[33]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[34]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[35]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[36]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[37]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFF47)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[38]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hF4F7FFFFF4F70000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[39]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h10D01FDF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h28E82BEB282BE8EB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_4_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_5_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEEEEEEEB22222228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_4 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_5 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[3]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFCF44CF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[40]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[41]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[42]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[43]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[44]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[45]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[46]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFCF44FFFFCF77)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[47]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[48]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[49]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88BB8B8B)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[4]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[50]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEB2228)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[51]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[52]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[53]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[54]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFEFFFFFFFEF0000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFF4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[55]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0407F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFF4FFF7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBFBFFF00BFBF00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[56]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[58]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair345" *) 
  LUT3 #(
    .INIT(8'h1D)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFBFBFFF00BFBF00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_3_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[57]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[59]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h88BB8B8B)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h1D1111111D11DDDD)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_2_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hEB2BFFFFFFFFFFFC)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_3_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[60]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h000001F1C0C001F1)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFEF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[61]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000200)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h02000020)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000001FF000001)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_4 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hFFFFFFEF)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h55555556)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h5555555555555556)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h56)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h5556)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0010FFFF00100000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_2_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_5_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_2_n_0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [63]),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00200000)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[63]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8B8B88BB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[14]_i_3_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[6]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8B888BBB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[15]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[7]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8BFF8B00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h7777777D44444441)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[16]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAFA0CFCFAFA0C0C0)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_4 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I1(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_7_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[8]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h04073437C4C7F4F7)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_1 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[11]_i_2_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[12]_i_2_n_0 ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[10]_i_2_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h8BFF8B00)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_9_n_0 ),
        .I2(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[13]_i_4_n_0 ),
        .I3(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[62]_i_8_n_0 ),
        .I4(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_3_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h22222228EEEEEEEB)) 
    \roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_3 
       (.I0(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[17]_i_4_n_0 ),
        .I1(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .I3(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .I4(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .I5(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[1]_i_4_n_0 ),
        .O(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_20_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_21_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_22_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_23_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_106 
       (.CI(\<const0>__0__0 ),
        .CO(roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_146_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_147_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_148_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_149_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111 
       (.CI(\<const0>__0__0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_150_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_151_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_152_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_153_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_31_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_32_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_33_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_34_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_19_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_36_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_37_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_38_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_39_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_1 ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_31_33 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_2_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_6_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_7_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_30_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_69_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_70_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_71_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_72_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_35_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_74_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_75_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_76_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_77_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_10_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_1 ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_21_29 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_4_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_11_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_12_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_13_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_5_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_14_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_15_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_16_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_17_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68 
       (.CI(roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[3]),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_68_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_107_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_108_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_109_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_110_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73 
       (.CI(\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_111_n_0 ),
        .CO({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_1 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_2 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg_reg[0]_i_73_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 ,\<const1>__0__0 }),
        .S({\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_112_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_113_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_114_n_0 ,\roundAndPackFloat64_shift64RightJammingexit_z0i_reg[0]_i_115_n_0 }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h0000FE02)) 
    roundAndPackFloat64_start_i_1
       (.I0(\main_inst/roundAndPackFloat64_start_reg_n_0 ),
        .I1(roundAndPackFloat64_start_i_2_n_0),
        .I2(\main_inst/roundAndPackFloat64_start ),
        .I3(roundAndPackFloat64_start_i_3_n_0),
        .I4(\main_inst/main_normalizeRoundAndPackFloat64exitii_214_reg ),
        .O(roundAndPackFloat64_start_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000200000080000)) 
    roundAndPackFloat64_start_i_2
       (.I0(roundAndPackFloat64_start_i_4_n_0),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\main_inst/cur_state_reg_n_0_[1] ),
        .I3(\main_inst/cur_state_reg_n_0_[3] ),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\main_inst/cur_state_reg_n_0_[6] ),
        .O(roundAndPackFloat64_start_i_2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFFFFFFFFDF)) 
    roundAndPackFloat64_start_i_3
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[1] ),
        .I5(\return_val[31]_i_3_n_0 ),
        .O(roundAndPackFloat64_start_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    roundAndPackFloat64_start_i_4
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .O(roundAndPackFloat64_start_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004000)) 
    roundAndPackFloat64_thread6_50_reg_i_1
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_10
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [36]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [37]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [34]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [35]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [39]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [38]),
        .O(roundAndPackFloat64_thread6_50_reg_i_10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_11
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [30]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [31]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [28]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [29]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [33]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [32]),
        .O(roundAndPackFloat64_thread6_50_reg_i_11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_12
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [18]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [19]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [16]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [17]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [21]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [20]),
        .O(roundAndPackFloat64_thread6_50_reg_i_12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_13
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [24]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [25]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [22]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [23]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [27]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [26]),
        .O(roundAndPackFloat64_thread6_50_reg_i_13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    roundAndPackFloat64_thread6_50_reg_i_14
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [4]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [5]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [6]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [7]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [8]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [9]),
        .O(roundAndPackFloat64_thread6_50_reg_i_14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    roundAndPackFloat64_thread6_50_reg_i_2
       (.I0(roundAndPackFloat64_thread6_50_reg_i_3_n_0),
        .I1(roundAndPackFloat64_thread6_50_reg_i_4_n_0),
        .I2(roundAndPackFloat64_thread6_50_reg_i_5_n_0),
        .I3(roundAndPackFloat64_thread6_50_reg_i_6_n_0),
        .I4(roundAndPackFloat64_thread6_50_reg_i_7_n_0),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_50 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_3
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [54]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [55]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [52]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [53]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [57]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [56]),
        .O(roundAndPackFloat64_thread6_50_reg_i_3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_4
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [60]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [61]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [58]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [59]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [63]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [62]),
        .O(roundAndPackFloat64_thread6_50_reg_i_4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_5
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [48]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [49]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [46]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [47]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [51]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [50]),
        .O(roundAndPackFloat64_thread6_50_reg_i_5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000100000000)) 
    roundAndPackFloat64_thread6_50_reg_i_6
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [14]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [15]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [13]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [12]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [11]),
        .I5(roundAndPackFloat64_thread6_50_reg_i_8_n_0),
        .O(roundAndPackFloat64_thread6_50_reg_i_6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h80000000)) 
    roundAndPackFloat64_thread6_50_reg_i_7
       (.I0(roundAndPackFloat64_thread6_50_reg_i_9_n_0),
        .I1(roundAndPackFloat64_thread6_50_reg_i_10_n_0),
        .I2(roundAndPackFloat64_thread6_50_reg_i_11_n_0),
        .I3(roundAndPackFloat64_thread6_50_reg_i_12_n_0),
        .I4(roundAndPackFloat64_thread6_50_reg_i_13_n_0),
        .O(roundAndPackFloat64_thread6_50_reg_i_7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00010000FFFFFFFF)) 
    roundAndPackFloat64_thread6_50_reg_i_8
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [1]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [0]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [3]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [2]),
        .I4(roundAndPackFloat64_thread6_50_reg_i_14_n_0),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43__0 ),
        .O(roundAndPackFloat64_thread6_50_reg_i_8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000001)) 
    roundAndPackFloat64_thread6_50_reg_i_9
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [42]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [43]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [40]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [41]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [45]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [44]),
        .O(roundAndPackFloat64_thread6_50_reg_i_9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \roundAndPackFloat64_thread6_55_reg[0]_i_1 
       (.I0(roundAndPackFloat64_thread6_55_reg),
        .I1(\roundAndPackFloat64_thread6_55_reg[0]_i_3_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_55 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0000FFFE0000)) 
    \roundAndPackFloat64_thread6_55_reg[0]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [0]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [3]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [4]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [2]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43__0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [1]),
        .O(roundAndPackFloat64_thread6_55_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF0000FFEF0000)) 
    \roundAndPackFloat64_thread6_55_reg[0]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [5]),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [8]),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [9]),
        .I3(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [7]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43__0 ),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_roundBits09_reg [6]),
        .O(\roundAndPackFloat64_thread6_55_reg[0]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \roundAndPackFloat64_thread6_55_reg[1]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[9] ),
        .O(\roundAndPackFloat64_thread6_55_reg[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[13]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_0 ),
        .CO(roundAndPackFloat64_thread6_55_reg_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [23:20]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[23] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[22] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[21] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[20] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[17]_i_1 
       (.CI(roundAndPackFloat64_thread6_55_reg_reg[3]),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [27:24]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[27] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[26] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[25] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[24] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[1]_i_1 
       (.CI(\<const0>__0__0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[9] ,\<const0>__0__0 }),
        .O({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [11],\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43__0 ,\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_6 ,\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_7 }),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[11] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_ ,\roundAndPackFloat64_thread6_55_reg[1]_i_4_n_0 ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[8] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[21]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[17]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [31:28]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[31] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[30] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[29] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[28] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[25]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[21]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [35:32]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[35] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[34] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[33] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[32] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[29]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[25]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [39:36]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[39] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[38] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[37] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[36] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[33]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[29]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [43:40]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[43] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[42] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[41] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[40] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[37]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[33]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [47:44]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[47] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[46] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[45] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[44] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[41]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[37]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [51:48]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[51] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[50] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[49] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[48] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[45]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[41]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [55:52]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[55] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[54] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[53] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[52] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[49]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[45]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [59:56]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[59] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[58] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[57] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[56] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[53]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[49]_i_1_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [63:60]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[63] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[62] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[61] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[60] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[5]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[1]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [15:12]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[15] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[14] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[13] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[12] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \roundAndPackFloat64_thread6_55_reg_reg[9]_i_1 
       (.CI(\roundAndPackFloat64_thread6_55_reg_reg[5]_i_1_n_0 ),
        .CO({\roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_0 ,\roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_1 ,\roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_2 ,\roundAndPackFloat64_thread6_55_reg_reg[9]_i_1_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_43 [19:16]),
        .S({\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[19] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[18] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[17] ,\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg_reg_n_0_[16] }));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0020000000000000)) 
    \roundAndPackFloat64_thread6_roundBits09_reg[9]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_35 ),
        .O(roundAndPackFloat64_thread6_roundBits09_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \roundAndPackFloat64_thread6_roundBits09_reg[9]_i_2 
       (.I0(roundAndPackFloat64_thread6_roundBits09_reg),
        .I1(\roundAndPackFloat64_thread6_roundBits09_reg[9]_i_3_n_0 ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000C00800)) 
    \roundAndPackFloat64_thread6_roundBits09_reg[9]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_39 ),
        .I1(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\roundAndPackFloat64_thread6_roundBits09_reg[9]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[10]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [10]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [10]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[11]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [11]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [11]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[12]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [12]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [12]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[13]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [13]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [13]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[14]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [14]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [14]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[15]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [15]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [15]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[16]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [16]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [16]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[17]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [17]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [17]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[18]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [18]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [18]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[19]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [19]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [19]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[20]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [20]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [20]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[21]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [21]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [21]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[22]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [22]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [22]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[23]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [23]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [23]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[24]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [24]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [24]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[25]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [25]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [25]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[26]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [26]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [26]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[27]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [27]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [27]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[28]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [28]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [28]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[29]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [29]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [29]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[30]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [30]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [30]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[31]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [31]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [31]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[32]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [32]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [32]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[33]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [33]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [33]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[34]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [34]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [34]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair354" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[35]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [35]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [35]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair353" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[36]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [36]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [36]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[37]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [37]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [37]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair351" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[38]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [38]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [38]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair347" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[39]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [39]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [39]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[40]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [40]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [40]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair357" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[41]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [41]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [41]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair346" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[42]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [42]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [42]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair344" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[43]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [43]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [43]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair356" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[44]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [44]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [44]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair343" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[45]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [45]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [45]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair342" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[46]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [46]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [46]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair341" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[47]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [47]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [47]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair340" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[48]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [48]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [48]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair339" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[49]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [49]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [49]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair336" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[50]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [50]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [50]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair335" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[51]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [51]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [51]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair334" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[52]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [52]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [52]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair333" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[53]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [53]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [53]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair355" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[54]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [54]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [54]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair332" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[55]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [55]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [55]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair328" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[56]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [56]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [56]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair352" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[57]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [57]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [57]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair326" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[58]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [58]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [58]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair350" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[59]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [59]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [59]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair349" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[60]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [60]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [60]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair348" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[61]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [61]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [61]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair325" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[62]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [62]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [62]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair323" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread6_zSig57_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [63]),
        .I1(roundAndPackFloat64_thread6_roundBits09_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5_reg [63]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread6_zSig57 [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[0]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_ ),
        .O(roundAndPackFloat64_thread_02_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000200)) 
    \roundAndPackFloat64_thread_02_reg[10]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I5(roundAndPackFloat64_thread_roundBits0_reg),
        .O(\roundAndPackFloat64_thread_02_reg[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[10]_i_2 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[10] ),
        .O(\roundAndPackFloat64_thread_02_reg[10]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000800000000)) 
    \roundAndPackFloat64_thread_02_reg[11]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\roundAndPackFloat64_thread_02_reg[11]_i_2_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I3(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[11] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'h0100)) 
    \roundAndPackFloat64_thread_02_reg[11]_i_2 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .O(\roundAndPackFloat64_thread_02_reg[11]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000080)) 
    \roundAndPackFloat64_thread_02_reg[11]_i_3 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_6_n_0 ),
        .I3(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ),
        .O(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFF000800000000)) 
    \roundAndPackFloat64_thread_02_reg[1]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\roundAndPackFloat64_thread_02_reg[11]_i_2_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I3(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I4(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I5(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[1] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_02 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[2]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[2] ),
        .O(\roundAndPackFloat64_thread_02_reg[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[3]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[3] ),
        .O(\roundAndPackFloat64_thread_02_reg[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[4]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[4] ),
        .O(\roundAndPackFloat64_thread_02_reg[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[5]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[5] ),
        .O(\roundAndPackFloat64_thread_02_reg[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[6]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[6] ),
        .O(\roundAndPackFloat64_thread_02_reg[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[7]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[7] ),
        .O(\roundAndPackFloat64_thread_02_reg[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[8]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[8] ),
        .O(\roundAndPackFloat64_thread_02_reg[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hF2)) 
    \roundAndPackFloat64_thread_02_reg[9]_i_1 
       (.I0(\roundAndPackFloat64_thread_02_reg[11]_i_3_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[9] ),
        .O(\roundAndPackFloat64_thread_02_reg[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[0]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_ ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_ ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_ ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [0]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[1]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[1] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[1] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[1] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [1]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[2]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[2] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[2] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[2] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [2]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[3]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[3] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[3] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[3] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [3]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[4]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[4] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[4] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[4] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [4]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[5]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[5] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[5] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[5] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [5]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[6]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[6] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[6] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[6] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [6]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[7]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[7] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[7] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[7] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [7]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[8]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[8] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[8] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF00040000)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_1 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I5(roundAndPackFloat64_thread_roundBits0_reg),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0_reg ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hB8BBB888)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_2 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_34_reg_reg_n_0_[9] ),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_1_reg_reg_n_0_[9] ),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_roundBits0 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hB)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_3 
       (.I0(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ),
        .I1(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ),
        .O(roundAndPackFloat64_thread_roundBits0_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000010000)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_4 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [3]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I2(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I3(\main_inst/roundAndPackFloat64/cur_state [1]),
        .I4(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I5(\main_inst/roundAndPackFloat64/roundAndPackFloat64_0_3 ),
        .O(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFCFFAFFFFFFFFFFF)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_5 
       (.I0(\main_inst/roundAndPackFloat64_arg_zExp_reg_n_0_[31] ),
        .I1(\main_inst/roundAndPackFloat64/roundAndPackFloat64_8_9 ),
        .I2(\main_inst/roundAndPackFloat64/cur_state [0]),
        .I3(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_6_n_0 ),
        .I4(\main_inst/roundAndPackFloat64/cur_state [4]),
        .I5(\main_inst/roundAndPackFloat64/cur_state [3]),
        .O(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h1)) 
    \roundAndPackFloat64_thread_roundBits0_reg[9]_i_6 
       (.I0(\main_inst/roundAndPackFloat64/cur_state [2]),
        .I1(\main_inst/roundAndPackFloat64/cur_state [1]),
        .O(\roundAndPackFloat64_thread_roundBits0_reg[9]_i_6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[10]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[10] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [10]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [10]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[11]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[11] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [11]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [11]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[12]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[12] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [12]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [12]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[13]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[13] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [13]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [13]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[14]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[14] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [14]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [14]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[15]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[15] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [15]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [15]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[16]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[16] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [16]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [16]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[17]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[17] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [17]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [17]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[18]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[18] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [18]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [18]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[19]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[19] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [19]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [19]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[20]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[20] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [20]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [20]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[21]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[21] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [21]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [21]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[22]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[22] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [22]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [22]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[23]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[23] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [23]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[24]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[24] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [24]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[25]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[25] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [25]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [25]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[26]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[26] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [26]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[27]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[27] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [27]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [27]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[28]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[28] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [28]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[29]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[29] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [29]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [29]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[30]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[30] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [30]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [30]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[31]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[31] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [31]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[32]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[32] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [32]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [32]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[33]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[33] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [33]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [33]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[34]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[34] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [34]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [34]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[35]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[35] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [35]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [35]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[36]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[36] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [36]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [36]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[37]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[37] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [37]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [37]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[38]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[38] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [38]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [38]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[39]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[39] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [39]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [39]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[40]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[40] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [40]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [40]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[41]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[41] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [41]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [41]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[42]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[42] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [42]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [42]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[43]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[43] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [43]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [43]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[44]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[44] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [44]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [44]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[45]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[45] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [45]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [45]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[46]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[46] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [46]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [46]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[47]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[47] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [47]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [47]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[48]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[48] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [48]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [48]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[49]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[49] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [49]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [49]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[50]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[50] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [50]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [50]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[51]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[51] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [51]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [51]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[52]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[52] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [52]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [52]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[53]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[53] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [53]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [53]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[54]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[54] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [54]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [54]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[55]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[55] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [55]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [55]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[56]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[56] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [56]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [56]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[57]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[57] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [57]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [57]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[58]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[58] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [58]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [58]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair324" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[59]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[59] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [59]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [59]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[60]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[60] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [60]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [60]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair337" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[61]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[61] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [61]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [61]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[62]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[62] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [62]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [62]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair338" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[63]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[63] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [63]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [63]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[8]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[8] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [8]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [8]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \roundAndPackFloat64_thread_zSig5_reg[9]_i_1 
       (.I0(\main_inst/roundAndPackFloat64_arg_zSig_reg_n_0_[9] ),
        .I1(roundAndPackFloat64_thread_roundBits0_reg),
        .I2(\main_inst/roundAndPackFloat64/roundAndPackFloat64_shift64RightJammingexit_z0i_reg [9]),
        .O(\main_inst/roundAndPackFloat64/roundAndPackFloat64_thread_zSig5 [9]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    \select_float_exception_flags_reg_a[1]_i_1 
       (.I0(\select_float_exception_flags_reg_a[1]_i_2_n_0 ),
        .I1(\select_float_exception_flags_reg_a[1]_i_3_n_0 ),
        .I2(\select_float_exception_flags_reg_a[1]_i_4_n_0 ),
        .I3(\select_float_exception_flags_reg_a[1]_i_5_n_0 ),
        .I4(memory_controller_address_a[23]),
        .O(\select_float_exception_flags_reg_a[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h40)) 
    \select_float_exception_flags_reg_a[1]_i_10 
       (.I0(\main_inst/cur_state_reg_n_0_[4] ),
        .I1(\main_inst/cur_state_reg_n_0_ ),
        .I2(\select_float_exception_flags_reg_a[1]_i_21_n_0 ),
        .O(select_float_exception_flags_reg_a));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004F40)) 
    \select_float_exception_flags_reg_a[1]_i_11 
       (.I0(select_float_exception_flags_reg_a),
        .I1(\main_inst/data2 [31]),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/main_1_scevgep_reg_reg_n_0_[31] ),
        .I4(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .O(memory_controller_address_a[31]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004F40)) 
    \select_float_exception_flags_reg_a[1]_i_13 
       (.I0(select_float_exception_flags_reg_a),
        .I1(\main_inst/data2 [26]),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/main_1_scevgep_reg_reg_n_0_[26] ),
        .I4(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .O(memory_controller_address_a[26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004F40)) 
    \select_float_exception_flags_reg_a[1]_i_14 
       (.I0(select_float_exception_flags_reg_a),
        .I1(\main_inst/data2 [28]),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/main_1_scevgep_reg_reg_n_0_[28] ),
        .I4(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .O(memory_controller_address_a[28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00FFE2FF00FFE200)) 
    \select_float_exception_flags_reg_a[1]_i_15 
       (.I0(\main_inst/data2 [24]),
        .I1(select_float_exception_flags_reg_a),
        .I2(\main_inst/roundAndPackFloat64_memory_controller_enable_a ),
        .I3(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I4(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .I5(\main_inst/main_1_scevgep_reg_reg_n_0_[24] ),
        .O(memory_controller_address_a[24]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000004000010081)) 
    \select_float_exception_flags_reg_a[1]_i_17 
       (.I0(\main_inst/cur_state_reg ),
        .I1(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I2(\main_inst/cur_state_reg_n_0_[3] ),
        .I3(\main_inst/cur_state_reg_n_0_[4] ),
        .I4(\main_inst/cur_state_reg_n_0_[5] ),
        .I5(\main_inst/cur_state_reg_n_0_[2] ),
        .O(\select_float_exception_flags_reg_a[1]_i_17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h000022A2)) 
    \select_float_exception_flags_reg_a[1]_i_18 
       (.I0(\main_inst/cur_state_reg_n_0_[3] ),
        .I1(\main_inst/cur_state_reg ),
        .I2(\main_inst/cur_state_reg_n_0_ ),
        .I3(\main_inst/cur_state_reg_n_0_[2] ),
        .I4(\main_inst/cur_state_reg_n_0_[4] ),
        .O(\select_float_exception_flags_reg_a[1]_i_18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF04045404)) 
    \select_float_exception_flags_reg_a[1]_i_2 
       (.I0(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .I1(\main_inst/main_1_scevgep_reg_reg_n_0_[30] ),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/data2 [30]),
        .I4(select_float_exception_flags_reg_a),
        .I5(memory_controller_address_a[31]),
        .O(\select_float_exception_flags_reg_a[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00480D00)) 
    \select_float_exception_flags_reg_a[1]_i_21 
       (.I0(\main_inst/cur_state_reg ),
        .I1(\main_inst/cur_state_reg_n_0_[3] ),
        .I2(\main_inst/cur_state_reg_n_0_[2] ),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .O(\select_float_exception_flags_reg_a[1]_i_21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \select_float_exception_flags_reg_a[1]_i_27 
       (.I0(\main_inst/main_1_scevgep_reg1 [24]),
        .O(\select_float_exception_flags_reg_a[1]_i_27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \select_float_exception_flags_reg_a[1]_i_28 
       (.I0(\main_inst/main_1_scevgep_reg1 [23]),
        .O(\select_float_exception_flags_reg_a[1]_i_28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF04045404)) 
    \select_float_exception_flags_reg_a[1]_i_3 
       (.I0(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .I1(\main_inst/main_1_scevgep_reg_reg_n_0_[27] ),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/data2 [27]),
        .I4(select_float_exception_flags_reg_a),
        .I5(memory_controller_address_a[26]),
        .O(\select_float_exception_flags_reg_a[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hFFFFFFFF04045404)) 
    \select_float_exception_flags_reg_a[1]_i_4 
       (.I0(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .I1(\main_inst/main_1_scevgep_reg_reg_n_0_[29] ),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/data2 [29]),
        .I4(select_float_exception_flags_reg_a),
        .I5(memory_controller_address_a[28]),
        .O(\select_float_exception_flags_reg_a[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'hAAA0A202AAAAA202)) 
    \select_float_exception_flags_reg_a[1]_i_5 
       (.I0(memory_controller_address_a[24]),
        .I1(\main_inst/main_1_scevgep_reg_reg_n_0_[25] ),
        .I2(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .I3(select_float_exception_flags_reg_a),
        .I4(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I5(\main_inst/data2 [25]),
        .O(\select_float_exception_flags_reg_a[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00004F40)) 
    \select_float_exception_flags_reg_a[1]_i_6 
       (.I0(select_float_exception_flags_reg_a),
        .I1(\main_inst/data2 [23]),
        .I2(\select_float_exception_flags_reg_a[1]_i_8_n_0 ),
        .I3(\main_inst/main_1_scevgep_reg_reg_n_0_ ),
        .I4(\select_float_exception_flags_reg_a[1]_i_7_n_0 ),
        .O(memory_controller_address_a[23]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h7)) 
    \select_float_exception_flags_reg_a[1]_i_7 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\select_float_exception_flags_reg_a[1]_i_17_n_0 ),
        .O(\select_float_exception_flags_reg_a[1]_i_7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hF6DFFFFF)) 
    \select_float_exception_flags_reg_a[1]_i_8 
       (.I0(\main_inst/cur_state_reg_n_0_ ),
        .I1(\main_inst/cur_state_reg_n_0_[2] ),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\main_inst/cur_state_reg[6]_rep_n_0 ),
        .I4(\select_float_exception_flags_reg_a[1]_i_18_n_0 ),
        .O(\select_float_exception_flags_reg_a[1]_i_8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \select_float_exception_flags_reg_a_reg[1]_i_12 
       (.CI(\select_float_exception_flags_reg_a_reg[1]_i_16_n_0 ),
        .CO(select_float_exception_flags_reg_a_reg),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(\main_inst/data2 [29:26]),
        .S(\main_inst/main_1_scevgep_reg1 [29:26]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \select_float_exception_flags_reg_a_reg[1]_i_16 
       (.CI(\<const0>__0__0 ),
        .CO({\select_float_exception_flags_reg_a_reg[1]_i_16_n_0 ,\select_float_exception_flags_reg_a_reg[1]_i_16_n_1 ,\select_float_exception_flags_reg_a_reg[1]_i_16_n_2 ,\select_float_exception_flags_reg_a_reg[1]_i_16_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\main_inst/main_1_scevgep_reg1 [24:23],\<const0>__0__0 }),
        .O({\main_inst/data2 [25:23],\select_float_exception_flags_reg_a_reg[1]_i_16_n_7 }),
        .S({\main_inst/main_1_scevgep_reg1 [25],\select_float_exception_flags_reg_a[1]_i_27_n_0 ,\select_float_exception_flags_reg_a[1]_i_28_n_0 ,\main_inst/main_1_scevgep_reg1 [22]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \select_float_exception_flags_reg_a_reg[1]_i_9 
       (.CI(select_float_exception_flags_reg_a_reg[3]),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O({\select_float_exception_flags_reg_a_reg[1]_i_9_n_4 ,\select_float_exception_flags_reg_a_reg[1]_i_9_n_5 ,\main_inst/data2 [31:30]}),
        .S({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_1_scevgep_reg1 [31:30]}));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00000100)) 
    \select_float_exception_flags_reg_b[1]_i_1 
       (.I0(\select_float_exception_flags_reg_b[1]_i_2_n_0 ),
        .I1(\select_float_exception_flags_reg_b[1]_i_3_n_0 ),
        .I2(\select_float_exception_flags_reg_b[1]_i_4_n_0 ),
        .I3(\select_float_exception_flags_reg_b[1]_i_5_n_0 ),
        .I4(memory_controller_address_b),
        .O(\select_float_exception_flags_reg_b[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \select_float_exception_flags_reg_b[1]_i_15 
       (.I0(\main_inst/main_1_scevgep_reg1 [25]),
        .O(select_float_exception_flags_reg_b));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000C0800000000)) 
    \select_float_exception_flags_reg_b[1]_i_2 
       (.I0(select_float_exception_flags_reg_b_reg[2]),
        .I1(memory_controller_enable_reg_b_i_2_n_0),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(select_float_exception_flags_reg_b_reg[3]),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(ram_reg_i_61_n_0),
        .O(\select_float_exception_flags_reg_b[1]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000C0800000000)) 
    \select_float_exception_flags_reg_b[1]_i_3 
       (.I0(\select_float_exception_flags_reg_b_reg[1]_i_8_n_4 ),
        .I1(memory_controller_enable_reg_b_i_2_n_0),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\select_float_exception_flags_reg_b_reg[1]_i_8_n_5 ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(ram_reg_i_61_n_0),
        .O(\select_float_exception_flags_reg_b[1]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000C0800000000)) 
    \select_float_exception_flags_reg_b[1]_i_4 
       (.I0(select_float_exception_flags_reg_b_reg[1]),
        .I1(memory_controller_enable_reg_b_i_2_n_0),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(select_float_exception_flags_reg_b_reg[0]),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(ram_reg_i_61_n_0),
        .O(\select_float_exception_flags_reg_b[1]_i_4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000800000000)) 
    \select_float_exception_flags_reg_b[1]_i_5 
       (.I0(\select_float_exception_flags_reg_b_reg[1]_i_8_n_7 ),
        .I1(memory_controller_enable_reg_b_i_2_n_0),
        .I2(\main_inst/cur_state_reg_n_0_[5] ),
        .I3(\select_float_exception_flags_reg_b_reg[1]_i_8_n_6 ),
        .I4(\main_inst/cur_state_reg_n_0_[6] ),
        .I5(ram_reg_i_61_n_0),
        .O(\select_float_exception_flags_reg_b[1]_i_5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h0000000000000020)) 
    \select_float_exception_flags_reg_b[1]_i_6 
       (.I0(ram_reg_i_61_n_0),
        .I1(\main_inst/cur_state_reg_n_0_[6] ),
        .I2(\main_inst/main_1_scevgep_reg1 [23]),
        .I3(\main_inst/cur_state_reg_n_0_[5] ),
        .I4(\main_inst/cur_state_reg ),
        .I5(\main_inst/cur_state_reg_n_0_[3] ),
        .O(memory_controller_address_b));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \select_float_exception_flags_reg_b_reg[1]_i_7 
       (.CI(\select_float_exception_flags_reg_b_reg[1]_i_8_n_0 ),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 ,\<const0>__0__0 }),
        .O(select_float_exception_flags_reg_b_reg),
        .S(\main_inst/main_1_scevgep_reg1 [31:28]));
  (* BOX_TYPE = "PRIMITIVE" *) 
  CARRY4 \select_float_exception_flags_reg_b_reg[1]_i_8 
       (.CI(\<const0>__0__0 ),
        .CO({\select_float_exception_flags_reg_b_reg[1]_i_8_n_0 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_1 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_2 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_3 }),
        .CYINIT(\<const0>__0__0 ),
        .DI({\<const0>__0__0 ,\<const0>__0__0 ,\main_inst/main_1_scevgep_reg1 [25],\<const0>__0__0 }),
        .O({\select_float_exception_flags_reg_b_reg[1]_i_8_n_4 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_5 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_6 ,\select_float_exception_flags_reg_b_reg[1]_i_8_n_7 }),
        .S({\main_inst/main_1_scevgep_reg1 [27:26],select_float_exception_flags_reg_b,\main_inst/main_1_scevgep_reg1 [24]}));
endmodule
