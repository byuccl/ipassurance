module bubblesort
   (clk,
    rst,
    load_i,
    writedata_i,
    readdata_o,
    start_i,
    done_o,
    interrupt_o,
    abort_i);
  input clk;
  input rst;
  input [48:0]load_i;
  input [391:0]writedata_i;
  output [391:0]readdata_o;
  input start_i;
  output done_o;
  output interrupt_o;
  input abort_i;

  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const0>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \<const1>__0__0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire STAGEN;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[0].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[10].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[11].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[12].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[13].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[14].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[15].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[16].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[17].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[18].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[19].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[1].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[1].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[1].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[1].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[1].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[20].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[21].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[22].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[23].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[24].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[25].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[26].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[27].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[28].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[29].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[2].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[30].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[31].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[32].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[33].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[34].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[35].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[36].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[37].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[38].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[39].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[3].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[40].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[41].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[42].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[43].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[44].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[45].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[46].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[47].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[48].stage/split_module/r_swap_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[4].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[5].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[6].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[7].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[8].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/p_0_in ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/p_1_out ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_bit1 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_bit2 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_compare_result ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_freeze_compare_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_run_reg_n_0_[0] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \STAGEN[9].stage/split_module/r_small_bit_reg_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire clk;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire done_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_pulses_reg_n_0_ ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_pulses_reg_n_0_[1] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_pulses_reg_n_0_[2] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_pulses_reg_n_0_[3] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_pulses_reg_n_0_[4] ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_run_delay ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \interrupt_module/r_swap_delay ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire interrupt_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [48:0]load_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [11:0]p_2_in;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_compare_result_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_count;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_data;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[0]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[1]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__0_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__10_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__11_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__12_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__13_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__14_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__15_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__16_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__17_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__18_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__19_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__20_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__21_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__22_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__23_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__24_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__25_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__26_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__27_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__28_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__29_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__30_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__31_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__32_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__33_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__34_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__35_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__36_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__37_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__38_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__39_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__40_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__41_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__42_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__43_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__44_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__45_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__46_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__47_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__4_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__5_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__6_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__7_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__8_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2__9_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_data[7]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_done_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_freeze_compare_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_job_done_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_large_bit_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_pulses;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_pulses0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[2]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[3]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[5]_i_2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_pulses[5]_i_3_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_run_late_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_run_late_66__0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__0_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__10_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__11_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__12_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__13_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__14_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__15_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__16_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__17_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__18_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__19_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__20_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__21_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__22_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__23_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__24_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__25_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__26_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__27_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__28_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__29_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__2_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__30_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__31_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__32_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__33_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__34_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__35_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__36_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__37_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__38_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__39_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__3_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__40_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__41_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__42_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__43_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__44_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__45_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__46_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__4_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__5_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__6_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__7_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__8_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1__9_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_small_bit_i_1_n_0;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_value_66;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire r_value_66_reg;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \r_value_66_reg[0]_srl2_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [391:0]readdata_o;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire rst;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[10]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[11]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[4]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[5]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[6]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[7]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[8]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_count[9]_i_1_n_0 ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire \run_module/r_job_done ;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire start_i;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_15;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_17;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_19;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_24;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_25;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_26;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_27;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_28;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_29;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_34;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_35;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_36;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_37;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_38;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_39;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_40;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_41;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_42;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_43;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_44;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_45;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_46;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_47;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_bit_up_9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_1;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_15;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_17;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_19;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_24;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_25;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_26;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_27;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_28;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_29;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_34;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_35;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_36;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_37;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_38;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_39;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_40;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_41;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_42;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_43;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_44;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_45;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_46;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_47;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_49;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_run_up_9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_10;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_11;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_12;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_13;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_14;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_15;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_16;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_17;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_18;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_19;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_2;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_20;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_21;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_22;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_23;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_24;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_25;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_26;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_27;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_28;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_29;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_3;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_30;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_31;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_32;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_33;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_34;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_35;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_36;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_37;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_38;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_39;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_4;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_40;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_41;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_42;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_43;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_44;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_45;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_46;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_47;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_48;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_5;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_6;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_7;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_8;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire w_swap_up_9;
  (* RTL_KEEP = "yes" *) (* STRUCTURAL_NETLIST = "yes" *) wire [391:0]writedata_i;

  (* BOX_TYPE = "PRIMITIVE" *) 
  GND GND
       (.G(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[0]_i_1_n_0 ),
        .Q(readdata_o[0]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[1]_i_1_n_0 ),
        .Q(readdata_o[1]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[2]_i_1_n_0 ),
        .Q(readdata_o[2]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[3]_i_1_n_0 ),
        .Q(readdata_o[3]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[4]_i_1_n_0 ),
        .Q(readdata_o[4]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[5]_i_1_n_0 ),
        .Q(readdata_o[5]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[6]_i_1_n_0 ),
        .Q(readdata_o[6]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1_n_0 ),
        .D(\r_data[7]_i_2_n_0 ),
        .Q(readdata_o[7]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[7]),
        .Q(STAGEN),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(STAGEN),
        .Q(w_bit_up_1),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run),
        .Q(\STAGEN[0].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[0].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[0].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_1),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[0]_i_1__9_n_0 ),
        .Q(readdata_o[80]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[1]_i_1__9_n_0 ),
        .Q(readdata_o[81]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[2]_i_1__9_n_0 ),
        .Q(readdata_o[82]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[3]_i_1__9_n_0 ),
        .Q(readdata_o[83]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[4]_i_1__9_n_0 ),
        .Q(readdata_o[84]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[5]_i_1__9_n_0 ),
        .Q(readdata_o[85]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[6]_i_1__9_n_0 ),
        .Q(readdata_o[86]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__9_n_0 ),
        .D(\r_data[7]_i_2__9_n_0 ),
        .Q(readdata_o[87]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_10),
        .Q(\STAGEN[10].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[87]),
        .Q(\STAGEN[10].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__8_n_0),
        .Q(\STAGEN[10].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__8_n_0),
        .Q(\STAGEN[10].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__8_n_0),
        .Q(w_bit_up_11),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_10),
        .Q(\STAGEN[10].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[10].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_11),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__8_n_0),
        .Q(\STAGEN[10].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_10),
        .Q(\STAGEN[10].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[10].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[10].stage/split_module/p_1_out ),
        .Q(w_swap_up_11),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[0]_i_1__10_n_0 ),
        .Q(readdata_o[88]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[1]_i_1__10_n_0 ),
        .Q(readdata_o[89]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[2]_i_1__10_n_0 ),
        .Q(readdata_o[90]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[3]_i_1__10_n_0 ),
        .Q(readdata_o[91]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[4]_i_1__10_n_0 ),
        .Q(readdata_o[92]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[5]_i_1__10_n_0 ),
        .Q(readdata_o[93]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[6]_i_1__10_n_0 ),
        .Q(readdata_o[94]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__10_n_0 ),
        .D(\r_data[7]_i_2__10_n_0 ),
        .Q(readdata_o[95]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_11),
        .Q(\STAGEN[11].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[95]),
        .Q(\STAGEN[11].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__9_n_0),
        .Q(\STAGEN[11].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__9_n_0),
        .Q(\STAGEN[11].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__9_n_0),
        .Q(w_bit_up_12),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_11),
        .Q(\STAGEN[11].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[11].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_12),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__9_n_0),
        .Q(\STAGEN[11].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_11),
        .Q(\STAGEN[11].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[11].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[11].stage/split_module/p_1_out ),
        .Q(w_swap_up_12),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[0]_i_1__11_n_0 ),
        .Q(readdata_o[96]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[1]_i_1__11_n_0 ),
        .Q(readdata_o[97]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[2]_i_1__11_n_0 ),
        .Q(readdata_o[98]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[3]_i_1__11_n_0 ),
        .Q(readdata_o[99]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[4]_i_1__11_n_0 ),
        .Q(readdata_o[100]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[5]_i_1__11_n_0 ),
        .Q(readdata_o[101]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[6]_i_1__11_n_0 ),
        .Q(readdata_o[102]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__11_n_0 ),
        .D(\r_data[7]_i_2__11_n_0 ),
        .Q(readdata_o[103]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_12),
        .Q(\STAGEN[12].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[103]),
        .Q(\STAGEN[12].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__10_n_0),
        .Q(\STAGEN[12].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__10_n_0),
        .Q(\STAGEN[12].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__10_n_0),
        .Q(w_bit_up_13),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_12),
        .Q(\STAGEN[12].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[12].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_13),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__10_n_0),
        .Q(\STAGEN[12].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_12),
        .Q(\STAGEN[12].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[12].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[12].stage/split_module/p_1_out ),
        .Q(w_swap_up_13),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[0]_i_1__12_n_0 ),
        .Q(readdata_o[104]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[1]_i_1__12_n_0 ),
        .Q(readdata_o[105]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[2]_i_1__12_n_0 ),
        .Q(readdata_o[106]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[3]_i_1__12_n_0 ),
        .Q(readdata_o[107]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[4]_i_1__12_n_0 ),
        .Q(readdata_o[108]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[5]_i_1__12_n_0 ),
        .Q(readdata_o[109]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[6]_i_1__12_n_0 ),
        .Q(readdata_o[110]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__12_n_0 ),
        .D(\r_data[7]_i_2__12_n_0 ),
        .Q(readdata_o[111]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_13),
        .Q(\STAGEN[13].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[111]),
        .Q(\STAGEN[13].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__11_n_0),
        .Q(\STAGEN[13].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__11_n_0),
        .Q(\STAGEN[13].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__11_n_0),
        .Q(w_bit_up_14),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_13),
        .Q(\STAGEN[13].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[13].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_14),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__11_n_0),
        .Q(\STAGEN[13].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_13),
        .Q(\STAGEN[13].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[13].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[13].stage/split_module/p_1_out ),
        .Q(w_swap_up_14),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[0]_i_1__13_n_0 ),
        .Q(readdata_o[112]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[1]_i_1__13_n_0 ),
        .Q(readdata_o[113]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[2]_i_1__13_n_0 ),
        .Q(readdata_o[114]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[3]_i_1__13_n_0 ),
        .Q(readdata_o[115]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[4]_i_1__13_n_0 ),
        .Q(readdata_o[116]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[5]_i_1__13_n_0 ),
        .Q(readdata_o[117]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[6]_i_1__13_n_0 ),
        .Q(readdata_o[118]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__13_n_0 ),
        .D(\r_data[7]_i_2__13_n_0 ),
        .Q(readdata_o[119]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_14),
        .Q(\STAGEN[14].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[119]),
        .Q(\STAGEN[14].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__12_n_0),
        .Q(\STAGEN[14].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__12_n_0),
        .Q(\STAGEN[14].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__12_n_0),
        .Q(w_bit_up_15),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_14),
        .Q(\STAGEN[14].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[14].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_15),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__12_n_0),
        .Q(\STAGEN[14].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_14),
        .Q(\STAGEN[14].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[14].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[14].stage/split_module/p_1_out ),
        .Q(w_swap_up_15),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[0]_i_1__14_n_0 ),
        .Q(readdata_o[120]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[1]_i_1__14_n_0 ),
        .Q(readdata_o[121]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[2]_i_1__14_n_0 ),
        .Q(readdata_o[122]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[3]_i_1__14_n_0 ),
        .Q(readdata_o[123]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[4]_i_1__14_n_0 ),
        .Q(readdata_o[124]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[5]_i_1__14_n_0 ),
        .Q(readdata_o[125]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[6]_i_1__14_n_0 ),
        .Q(readdata_o[126]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__14_n_0 ),
        .D(\r_data[7]_i_2__14_n_0 ),
        .Q(readdata_o[127]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_15),
        .Q(\STAGEN[15].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[127]),
        .Q(\STAGEN[15].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__13_n_0),
        .Q(\STAGEN[15].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__13_n_0),
        .Q(\STAGEN[15].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__13_n_0),
        .Q(w_bit_up_16),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_15),
        .Q(\STAGEN[15].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[15].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_16),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__13_n_0),
        .Q(\STAGEN[15].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_15),
        .Q(\STAGEN[15].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[15].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[15].stage/split_module/p_1_out ),
        .Q(w_swap_up_16),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[0]_i_1__15_n_0 ),
        .Q(readdata_o[128]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[1]_i_1__15_n_0 ),
        .Q(readdata_o[129]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[2]_i_1__15_n_0 ),
        .Q(readdata_o[130]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[3]_i_1__15_n_0 ),
        .Q(readdata_o[131]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[4]_i_1__15_n_0 ),
        .Q(readdata_o[132]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[5]_i_1__15_n_0 ),
        .Q(readdata_o[133]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[6]_i_1__15_n_0 ),
        .Q(readdata_o[134]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__15_n_0 ),
        .D(\r_data[7]_i_2__15_n_0 ),
        .Q(readdata_o[135]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_16),
        .Q(\STAGEN[16].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[135]),
        .Q(\STAGEN[16].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__14_n_0),
        .Q(\STAGEN[16].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__14_n_0),
        .Q(\STAGEN[16].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__14_n_0),
        .Q(w_bit_up_17),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_16),
        .Q(\STAGEN[16].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[16].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_17),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__14_n_0),
        .Q(\STAGEN[16].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_16),
        .Q(\STAGEN[16].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[16].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[16].stage/split_module/p_1_out ),
        .Q(w_swap_up_17),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[0]_i_1__16_n_0 ),
        .Q(readdata_o[136]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[1]_i_1__16_n_0 ),
        .Q(readdata_o[137]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[2]_i_1__16_n_0 ),
        .Q(readdata_o[138]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[3]_i_1__16_n_0 ),
        .Q(readdata_o[139]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[4]_i_1__16_n_0 ),
        .Q(readdata_o[140]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[5]_i_1__16_n_0 ),
        .Q(readdata_o[141]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[6]_i_1__16_n_0 ),
        .Q(readdata_o[142]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__16_n_0 ),
        .D(\r_data[7]_i_2__16_n_0 ),
        .Q(readdata_o[143]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_17),
        .Q(\STAGEN[17].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[143]),
        .Q(\STAGEN[17].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__15_n_0),
        .Q(\STAGEN[17].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__15_n_0),
        .Q(\STAGEN[17].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__15_n_0),
        .Q(w_bit_up_18),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_17),
        .Q(\STAGEN[17].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[17].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_18),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__15_n_0),
        .Q(\STAGEN[17].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_17),
        .Q(\STAGEN[17].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[17].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[17].stage/split_module/p_1_out ),
        .Q(w_swap_up_18),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[0]_i_1__17_n_0 ),
        .Q(readdata_o[144]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[1]_i_1__17_n_0 ),
        .Q(readdata_o[145]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[2]_i_1__17_n_0 ),
        .Q(readdata_o[146]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[3]_i_1__17_n_0 ),
        .Q(readdata_o[147]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[4]_i_1__17_n_0 ),
        .Q(readdata_o[148]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[5]_i_1__17_n_0 ),
        .Q(readdata_o[149]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[6]_i_1__17_n_0 ),
        .Q(readdata_o[150]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__17_n_0 ),
        .D(\r_data[7]_i_2__17_n_0 ),
        .Q(readdata_o[151]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_18),
        .Q(\STAGEN[18].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[151]),
        .Q(\STAGEN[18].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__16_n_0),
        .Q(\STAGEN[18].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__16_n_0),
        .Q(\STAGEN[18].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__16_n_0),
        .Q(w_bit_up_19),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_18),
        .Q(\STAGEN[18].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[18].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_19),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__16_n_0),
        .Q(\STAGEN[18].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_18),
        .Q(\STAGEN[18].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[18].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[18].stage/split_module/p_1_out ),
        .Q(w_swap_up_19),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[0]_i_1__18_n_0 ),
        .Q(readdata_o[152]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[1]_i_1__18_n_0 ),
        .Q(readdata_o[153]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[2]_i_1__18_n_0 ),
        .Q(readdata_o[154]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[3]_i_1__18_n_0 ),
        .Q(readdata_o[155]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[4]_i_1__18_n_0 ),
        .Q(readdata_o[156]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[5]_i_1__18_n_0 ),
        .Q(readdata_o[157]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[6]_i_1__18_n_0 ),
        .Q(readdata_o[158]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__18_n_0 ),
        .D(\r_data[7]_i_2__18_n_0 ),
        .Q(readdata_o[159]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_19),
        .Q(\STAGEN[19].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[159]),
        .Q(\STAGEN[19].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__17_n_0),
        .Q(\STAGEN[19].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__17_n_0),
        .Q(\STAGEN[19].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__17_n_0),
        .Q(w_bit_up_20),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_19),
        .Q(\STAGEN[19].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[19].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_20),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__17_n_0),
        .Q(\STAGEN[19].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_19),
        .Q(\STAGEN[19].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[19].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[19].stage/split_module/p_1_out ),
        .Q(w_swap_up_20),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(r_data),
        .Q(readdata_o[8]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[1]_i_1__0_n_0 ),
        .Q(readdata_o[9]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[2]_i_1__0_n_0 ),
        .Q(readdata_o[10]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[3]_i_1__0_n_0 ),
        .Q(readdata_o[11]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[4]_i_1__0_n_0 ),
        .Q(readdata_o[12]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[5]_i_1__0_n_0 ),
        .Q(readdata_o[13]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[6]_i_1__0_n_0 ),
        .Q(readdata_o[14]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__0_n_0 ),
        .D(\r_data[7]_i_2__0_n_0 ),
        .Q(readdata_o[15]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_1),
        .Q(\STAGEN[1].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[15]),
        .Q(\STAGEN[1].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1_n_0),
        .Q(\STAGEN[1].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1_n_0),
        .Q(\STAGEN[1].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1_n_0),
        .Q(w_bit_up_2),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_1),
        .Q(\STAGEN[1].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[1].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_2),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1_n_0),
        .Q(r_small_bit),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[1].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[1].stage/split_module/r_compare_result ),
        .Q(w_swap_up_2),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[0]_i_1__19_n_0 ),
        .Q(readdata_o[160]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[1]_i_1__19_n_0 ),
        .Q(readdata_o[161]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[2]_i_1__19_n_0 ),
        .Q(readdata_o[162]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[3]_i_1__19_n_0 ),
        .Q(readdata_o[163]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[4]_i_1__19_n_0 ),
        .Q(readdata_o[164]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[5]_i_1__19_n_0 ),
        .Q(readdata_o[165]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[6]_i_1__19_n_0 ),
        .Q(readdata_o[166]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__19_n_0 ),
        .D(\r_data[7]_i_2__19_n_0 ),
        .Q(readdata_o[167]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_20),
        .Q(\STAGEN[20].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[167]),
        .Q(\STAGEN[20].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__18_n_0),
        .Q(\STAGEN[20].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__18_n_0),
        .Q(\STAGEN[20].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__18_n_0),
        .Q(w_bit_up_21),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_20),
        .Q(\STAGEN[20].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[20].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_21),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__18_n_0),
        .Q(\STAGEN[20].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_20),
        .Q(\STAGEN[20].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[20].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[20].stage/split_module/p_1_out ),
        .Q(w_swap_up_21),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[0]_i_1__20_n_0 ),
        .Q(readdata_o[168]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[1]_i_1__20_n_0 ),
        .Q(readdata_o[169]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[2]_i_1__20_n_0 ),
        .Q(readdata_o[170]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[3]_i_1__20_n_0 ),
        .Q(readdata_o[171]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[4]_i_1__20_n_0 ),
        .Q(readdata_o[172]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[5]_i_1__20_n_0 ),
        .Q(readdata_o[173]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[6]_i_1__20_n_0 ),
        .Q(readdata_o[174]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__20_n_0 ),
        .D(\r_data[7]_i_2__20_n_0 ),
        .Q(readdata_o[175]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_21),
        .Q(\STAGEN[21].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[175]),
        .Q(\STAGEN[21].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__19_n_0),
        .Q(\STAGEN[21].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__19_n_0),
        .Q(\STAGEN[21].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__19_n_0),
        .Q(w_bit_up_22),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_21),
        .Q(\STAGEN[21].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[21].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_22),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__19_n_0),
        .Q(\STAGEN[21].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_21),
        .Q(\STAGEN[21].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[21].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[21].stage/split_module/p_1_out ),
        .Q(w_swap_up_22),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[0]_i_1__21_n_0 ),
        .Q(readdata_o[176]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[1]_i_1__21_n_0 ),
        .Q(readdata_o[177]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[2]_i_1__21_n_0 ),
        .Q(readdata_o[178]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[3]_i_1__21_n_0 ),
        .Q(readdata_o[179]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[4]_i_1__21_n_0 ),
        .Q(readdata_o[180]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[5]_i_1__21_n_0 ),
        .Q(readdata_o[181]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[6]_i_1__21_n_0 ),
        .Q(readdata_o[182]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__21_n_0 ),
        .D(\r_data[7]_i_2__21_n_0 ),
        .Q(readdata_o[183]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_22),
        .Q(\STAGEN[22].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[183]),
        .Q(\STAGEN[22].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__20_n_0),
        .Q(\STAGEN[22].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__20_n_0),
        .Q(\STAGEN[22].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__20_n_0),
        .Q(w_bit_up_23),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_22),
        .Q(\STAGEN[22].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[22].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_23),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__20_n_0),
        .Q(\STAGEN[22].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_22),
        .Q(\STAGEN[22].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[22].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[22].stage/split_module/p_1_out ),
        .Q(w_swap_up_23),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[0]_i_1__22_n_0 ),
        .Q(readdata_o[184]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[1]_i_1__22_n_0 ),
        .Q(readdata_o[185]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[2]_i_1__22_n_0 ),
        .Q(readdata_o[186]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[3]_i_1__22_n_0 ),
        .Q(readdata_o[187]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[4]_i_1__22_n_0 ),
        .Q(readdata_o[188]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[5]_i_1__22_n_0 ),
        .Q(readdata_o[189]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[6]_i_1__22_n_0 ),
        .Q(readdata_o[190]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__22_n_0 ),
        .D(\r_data[7]_i_2__22_n_0 ),
        .Q(readdata_o[191]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_23),
        .Q(\STAGEN[23].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[191]),
        .Q(\STAGEN[23].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__21_n_0),
        .Q(\STAGEN[23].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__21_n_0),
        .Q(\STAGEN[23].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__21_n_0),
        .Q(w_bit_up_24),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_23),
        .Q(\STAGEN[23].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[23].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_24),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__21_n_0),
        .Q(\STAGEN[23].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_23),
        .Q(\STAGEN[23].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[23].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[23].stage/split_module/p_1_out ),
        .Q(w_swap_up_24),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[0]_i_1__23_n_0 ),
        .Q(readdata_o[192]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[1]_i_1__23_n_0 ),
        .Q(readdata_o[193]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[2]_i_1__23_n_0 ),
        .Q(readdata_o[194]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[3]_i_1__23_n_0 ),
        .Q(readdata_o[195]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[4]_i_1__23_n_0 ),
        .Q(readdata_o[196]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[5]_i_1__23_n_0 ),
        .Q(readdata_o[197]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[6]_i_1__23_n_0 ),
        .Q(readdata_o[198]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__23_n_0 ),
        .D(\r_data[7]_i_2__23_n_0 ),
        .Q(readdata_o[199]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_24),
        .Q(\STAGEN[24].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[199]),
        .Q(\STAGEN[24].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__22_n_0),
        .Q(\STAGEN[24].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__22_n_0),
        .Q(\STAGEN[24].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__22_n_0),
        .Q(w_bit_up_25),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_24),
        .Q(\STAGEN[24].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[24].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_25),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__22_n_0),
        .Q(\STAGEN[24].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_24),
        .Q(\STAGEN[24].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[24].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[24].stage/split_module/p_1_out ),
        .Q(w_swap_up_25),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[0]_i_1__24_n_0 ),
        .Q(readdata_o[200]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[1]_i_1__24_n_0 ),
        .Q(readdata_o[201]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[2]_i_1__24_n_0 ),
        .Q(readdata_o[202]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[3]_i_1__24_n_0 ),
        .Q(readdata_o[203]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[4]_i_1__24_n_0 ),
        .Q(readdata_o[204]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[5]_i_1__24_n_0 ),
        .Q(readdata_o[205]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[6]_i_1__24_n_0 ),
        .Q(readdata_o[206]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__24_n_0 ),
        .D(\r_data[7]_i_2__24_n_0 ),
        .Q(readdata_o[207]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_25),
        .Q(\STAGEN[25].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[207]),
        .Q(\STAGEN[25].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__23_n_0),
        .Q(\STAGEN[25].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__23_n_0),
        .Q(\STAGEN[25].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__23_n_0),
        .Q(w_bit_up_26),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_25),
        .Q(\STAGEN[25].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[25].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_26),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__23_n_0),
        .Q(\STAGEN[25].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_25),
        .Q(\STAGEN[25].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[25].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[25].stage/split_module/p_1_out ),
        .Q(w_swap_up_26),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[0]_i_1__25_n_0 ),
        .Q(readdata_o[208]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[1]_i_1__25_n_0 ),
        .Q(readdata_o[209]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[2]_i_1__25_n_0 ),
        .Q(readdata_o[210]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[3]_i_1__25_n_0 ),
        .Q(readdata_o[211]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[4]_i_1__25_n_0 ),
        .Q(readdata_o[212]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[5]_i_1__25_n_0 ),
        .Q(readdata_o[213]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[6]_i_1__25_n_0 ),
        .Q(readdata_o[214]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__25_n_0 ),
        .D(\r_data[7]_i_2__25_n_0 ),
        .Q(readdata_o[215]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_26),
        .Q(\STAGEN[26].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[215]),
        .Q(\STAGEN[26].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__24_n_0),
        .Q(\STAGEN[26].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__24_n_0),
        .Q(\STAGEN[26].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__24_n_0),
        .Q(w_bit_up_27),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_26),
        .Q(\STAGEN[26].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[26].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_27),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__24_n_0),
        .Q(\STAGEN[26].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_26),
        .Q(\STAGEN[26].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[26].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[26].stage/split_module/p_1_out ),
        .Q(w_swap_up_27),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[0]_i_1__26_n_0 ),
        .Q(readdata_o[216]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[1]_i_1__26_n_0 ),
        .Q(readdata_o[217]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[2]_i_1__26_n_0 ),
        .Q(readdata_o[218]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[3]_i_1__26_n_0 ),
        .Q(readdata_o[219]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[4]_i_1__26_n_0 ),
        .Q(readdata_o[220]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[5]_i_1__26_n_0 ),
        .Q(readdata_o[221]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[6]_i_1__26_n_0 ),
        .Q(readdata_o[222]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__26_n_0 ),
        .D(\r_data[7]_i_2__26_n_0 ),
        .Q(readdata_o[223]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_27),
        .Q(\STAGEN[27].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[223]),
        .Q(\STAGEN[27].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__25_n_0),
        .Q(\STAGEN[27].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__25_n_0),
        .Q(\STAGEN[27].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__25_n_0),
        .Q(w_bit_up_28),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_27),
        .Q(\STAGEN[27].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[27].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_28),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__25_n_0),
        .Q(\STAGEN[27].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_27),
        .Q(\STAGEN[27].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[27].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[27].stage/split_module/p_1_out ),
        .Q(w_swap_up_28),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[0]_i_1__27_n_0 ),
        .Q(readdata_o[224]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[1]_i_1__27_n_0 ),
        .Q(readdata_o[225]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[2]_i_1__27_n_0 ),
        .Q(readdata_o[226]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[3]_i_1__27_n_0 ),
        .Q(readdata_o[227]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[4]_i_1__27_n_0 ),
        .Q(readdata_o[228]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[5]_i_1__27_n_0 ),
        .Q(readdata_o[229]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[6]_i_1__27_n_0 ),
        .Q(readdata_o[230]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__27_n_0 ),
        .D(\r_data[7]_i_2__27_n_0 ),
        .Q(readdata_o[231]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_28),
        .Q(\STAGEN[28].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[231]),
        .Q(\STAGEN[28].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__26_n_0),
        .Q(\STAGEN[28].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__26_n_0),
        .Q(\STAGEN[28].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__26_n_0),
        .Q(w_bit_up_29),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_28),
        .Q(\STAGEN[28].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[28].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_29),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__26_n_0),
        .Q(\STAGEN[28].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_28),
        .Q(\STAGEN[28].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[28].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[28].stage/split_module/p_1_out ),
        .Q(w_swap_up_29),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[0]_i_1__28_n_0 ),
        .Q(readdata_o[232]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[1]_i_1__28_n_0 ),
        .Q(readdata_o[233]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[2]_i_1__28_n_0 ),
        .Q(readdata_o[234]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[3]_i_1__28_n_0 ),
        .Q(readdata_o[235]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[4]_i_1__28_n_0 ),
        .Q(readdata_o[236]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[5]_i_1__28_n_0 ),
        .Q(readdata_o[237]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[6]_i_1__28_n_0 ),
        .Q(readdata_o[238]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__28_n_0 ),
        .D(\r_data[7]_i_2__28_n_0 ),
        .Q(readdata_o[239]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_29),
        .Q(\STAGEN[29].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[239]),
        .Q(\STAGEN[29].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__27_n_0),
        .Q(\STAGEN[29].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__27_n_0),
        .Q(\STAGEN[29].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__27_n_0),
        .Q(w_bit_up_30),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_29),
        .Q(\STAGEN[29].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[29].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_30),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__27_n_0),
        .Q(\STAGEN[29].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_29),
        .Q(\STAGEN[29].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[29].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[29].stage/split_module/p_1_out ),
        .Q(w_swap_up_30),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[0]_i_1__1_n_0 ),
        .Q(readdata_o[16]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[1]_i_1__1_n_0 ),
        .Q(readdata_o[17]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[2]_i_1__1_n_0 ),
        .Q(readdata_o[18]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[3]_i_1__1_n_0 ),
        .Q(readdata_o[19]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[4]_i_1__1_n_0 ),
        .Q(readdata_o[20]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[5]_i_1__1_n_0 ),
        .Q(readdata_o[21]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[6]_i_1__1_n_0 ),
        .Q(readdata_o[22]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__1_n_0 ),
        .D(\r_data[7]_i_2__1_n_0 ),
        .Q(readdata_o[23]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_2),
        .Q(\STAGEN[2].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[23]),
        .Q(\STAGEN[2].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__0_n_0),
        .Q(\STAGEN[2].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__0_n_0),
        .Q(\STAGEN[2].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__0_n_0),
        .Q(w_bit_up_3),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_2),
        .Q(\STAGEN[2].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[2].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_3),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__0_n_0),
        .Q(\STAGEN[2].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_2),
        .Q(\STAGEN[2].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[2].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[2].stage/split_module/p_1_out ),
        .Q(w_swap_up_3),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[0]_i_1__29_n_0 ),
        .Q(readdata_o[240]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[1]_i_1__29_n_0 ),
        .Q(readdata_o[241]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[2]_i_1__29_n_0 ),
        .Q(readdata_o[242]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[3]_i_1__29_n_0 ),
        .Q(readdata_o[243]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[4]_i_1__29_n_0 ),
        .Q(readdata_o[244]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[5]_i_1__29_n_0 ),
        .Q(readdata_o[245]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[6]_i_1__29_n_0 ),
        .Q(readdata_o[246]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__29_n_0 ),
        .D(\r_data[7]_i_2__29_n_0 ),
        .Q(readdata_o[247]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_30),
        .Q(\STAGEN[30].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[247]),
        .Q(\STAGEN[30].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__28_n_0),
        .Q(\STAGEN[30].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__28_n_0),
        .Q(\STAGEN[30].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__28_n_0),
        .Q(w_bit_up_31),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_30),
        .Q(\STAGEN[30].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[30].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_31),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__28_n_0),
        .Q(\STAGEN[30].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_30),
        .Q(\STAGEN[30].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[30].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[30].stage/split_module/p_1_out ),
        .Q(w_swap_up_31),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[0]_i_1__30_n_0 ),
        .Q(readdata_o[248]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[1]_i_1__30_n_0 ),
        .Q(readdata_o[249]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[2]_i_1__30_n_0 ),
        .Q(readdata_o[250]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[3]_i_1__30_n_0 ),
        .Q(readdata_o[251]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[4]_i_1__30_n_0 ),
        .Q(readdata_o[252]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[5]_i_1__30_n_0 ),
        .Q(readdata_o[253]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[6]_i_1__30_n_0 ),
        .Q(readdata_o[254]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__30_n_0 ),
        .D(\r_data[7]_i_2__30_n_0 ),
        .Q(readdata_o[255]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_31),
        .Q(\STAGEN[31].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[255]),
        .Q(\STAGEN[31].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__29_n_0),
        .Q(\STAGEN[31].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__29_n_0),
        .Q(\STAGEN[31].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__29_n_0),
        .Q(w_bit_up_32),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_31),
        .Q(\STAGEN[31].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[31].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_32),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__29_n_0),
        .Q(\STAGEN[31].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_31),
        .Q(\STAGEN[31].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[31].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[31].stage/split_module/p_1_out ),
        .Q(w_swap_up_32),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[0]_i_1__31_n_0 ),
        .Q(readdata_o[256]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[1]_i_1__31_n_0 ),
        .Q(readdata_o[257]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[2]_i_1__31_n_0 ),
        .Q(readdata_o[258]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[3]_i_1__31_n_0 ),
        .Q(readdata_o[259]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[4]_i_1__31_n_0 ),
        .Q(readdata_o[260]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[5]_i_1__31_n_0 ),
        .Q(readdata_o[261]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[6]_i_1__31_n_0 ),
        .Q(readdata_o[262]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__31_n_0 ),
        .D(\r_data[7]_i_2__31_n_0 ),
        .Q(readdata_o[263]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_32),
        .Q(\STAGEN[32].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[263]),
        .Q(\STAGEN[32].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__30_n_0),
        .Q(\STAGEN[32].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__30_n_0),
        .Q(\STAGEN[32].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__30_n_0),
        .Q(w_bit_up_33),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_32),
        .Q(\STAGEN[32].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[32].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_33),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__30_n_0),
        .Q(\STAGEN[32].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_32),
        .Q(\STAGEN[32].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[32].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[32].stage/split_module/p_1_out ),
        .Q(w_swap_up_33),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[0]_i_1__32_n_0 ),
        .Q(readdata_o[264]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[1]_i_1__32_n_0 ),
        .Q(readdata_o[265]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[2]_i_1__32_n_0 ),
        .Q(readdata_o[266]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[3]_i_1__32_n_0 ),
        .Q(readdata_o[267]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[4]_i_1__32_n_0 ),
        .Q(readdata_o[268]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[5]_i_1__32_n_0 ),
        .Q(readdata_o[269]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[6]_i_1__32_n_0 ),
        .Q(readdata_o[270]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__32_n_0 ),
        .D(\r_data[7]_i_2__32_n_0 ),
        .Q(readdata_o[271]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_33),
        .Q(\STAGEN[33].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[271]),
        .Q(\STAGEN[33].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__31_n_0),
        .Q(\STAGEN[33].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__31_n_0),
        .Q(\STAGEN[33].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__31_n_0),
        .Q(w_bit_up_34),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_33),
        .Q(\STAGEN[33].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[33].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_34),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__31_n_0),
        .Q(\STAGEN[33].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_33),
        .Q(\STAGEN[33].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[33].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[33].stage/split_module/p_1_out ),
        .Q(w_swap_up_34),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[0]_i_1__33_n_0 ),
        .Q(readdata_o[272]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[1]_i_1__33_n_0 ),
        .Q(readdata_o[273]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[2]_i_1__33_n_0 ),
        .Q(readdata_o[274]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[3]_i_1__33_n_0 ),
        .Q(readdata_o[275]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[4]_i_1__33_n_0 ),
        .Q(readdata_o[276]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[5]_i_1__33_n_0 ),
        .Q(readdata_o[277]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[6]_i_1__33_n_0 ),
        .Q(readdata_o[278]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__33_n_0 ),
        .D(\r_data[7]_i_2__33_n_0 ),
        .Q(readdata_o[279]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_34),
        .Q(\STAGEN[34].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[279]),
        .Q(\STAGEN[34].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__32_n_0),
        .Q(\STAGEN[34].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__32_n_0),
        .Q(\STAGEN[34].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__32_n_0),
        .Q(w_bit_up_35),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_34),
        .Q(\STAGEN[34].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[34].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_35),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__32_n_0),
        .Q(\STAGEN[34].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_34),
        .Q(\STAGEN[34].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[34].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[34].stage/split_module/p_1_out ),
        .Q(w_swap_up_35),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[0]_i_1__34_n_0 ),
        .Q(readdata_o[280]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[1]_i_1__34_n_0 ),
        .Q(readdata_o[281]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[2]_i_1__34_n_0 ),
        .Q(readdata_o[282]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[3]_i_1__34_n_0 ),
        .Q(readdata_o[283]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[4]_i_1__34_n_0 ),
        .Q(readdata_o[284]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[5]_i_1__34_n_0 ),
        .Q(readdata_o[285]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[6]_i_1__34_n_0 ),
        .Q(readdata_o[286]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__34_n_0 ),
        .D(\r_data[7]_i_2__34_n_0 ),
        .Q(readdata_o[287]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_35),
        .Q(\STAGEN[35].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[287]),
        .Q(\STAGEN[35].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__33_n_0),
        .Q(\STAGEN[35].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__33_n_0),
        .Q(\STAGEN[35].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__33_n_0),
        .Q(w_bit_up_36),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_35),
        .Q(\STAGEN[35].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[35].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_36),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__33_n_0),
        .Q(\STAGEN[35].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_35),
        .Q(\STAGEN[35].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[35].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[35].stage/split_module/p_1_out ),
        .Q(w_swap_up_36),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[0]_i_1__35_n_0 ),
        .Q(readdata_o[288]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[1]_i_1__35_n_0 ),
        .Q(readdata_o[289]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[2]_i_1__35_n_0 ),
        .Q(readdata_o[290]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[3]_i_1__35_n_0 ),
        .Q(readdata_o[291]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[4]_i_1__35_n_0 ),
        .Q(readdata_o[292]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[5]_i_1__35_n_0 ),
        .Q(readdata_o[293]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[6]_i_1__35_n_0 ),
        .Q(readdata_o[294]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__35_n_0 ),
        .D(\r_data[7]_i_2__35_n_0 ),
        .Q(readdata_o[295]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_36),
        .Q(\STAGEN[36].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[295]),
        .Q(\STAGEN[36].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__34_n_0),
        .Q(\STAGEN[36].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__34_n_0),
        .Q(\STAGEN[36].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__34_n_0),
        .Q(w_bit_up_37),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_36),
        .Q(\STAGEN[36].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[36].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_37),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__34_n_0),
        .Q(\STAGEN[36].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_36),
        .Q(\STAGEN[36].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[36].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[36].stage/split_module/p_1_out ),
        .Q(w_swap_up_37),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[0]_i_1__36_n_0 ),
        .Q(readdata_o[296]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[1]_i_1__36_n_0 ),
        .Q(readdata_o[297]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[2]_i_1__36_n_0 ),
        .Q(readdata_o[298]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[3]_i_1__36_n_0 ),
        .Q(readdata_o[299]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[4]_i_1__36_n_0 ),
        .Q(readdata_o[300]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[5]_i_1__36_n_0 ),
        .Q(readdata_o[301]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[6]_i_1__36_n_0 ),
        .Q(readdata_o[302]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__36_n_0 ),
        .D(\r_data[7]_i_2__36_n_0 ),
        .Q(readdata_o[303]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_37),
        .Q(\STAGEN[37].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[303]),
        .Q(\STAGEN[37].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__35_n_0),
        .Q(\STAGEN[37].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__35_n_0),
        .Q(\STAGEN[37].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__35_n_0),
        .Q(w_bit_up_38),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_37),
        .Q(\STAGEN[37].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[37].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_38),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__35_n_0),
        .Q(\STAGEN[37].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_37),
        .Q(\STAGEN[37].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[37].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[37].stage/split_module/p_1_out ),
        .Q(w_swap_up_38),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[0]_i_1__37_n_0 ),
        .Q(readdata_o[304]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[1]_i_1__37_n_0 ),
        .Q(readdata_o[305]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[2]_i_1__37_n_0 ),
        .Q(readdata_o[306]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[3]_i_1__37_n_0 ),
        .Q(readdata_o[307]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[4]_i_1__37_n_0 ),
        .Q(readdata_o[308]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[5]_i_1__37_n_0 ),
        .Q(readdata_o[309]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[6]_i_1__37_n_0 ),
        .Q(readdata_o[310]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__37_n_0 ),
        .D(\r_data[7]_i_2__37_n_0 ),
        .Q(readdata_o[311]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_38),
        .Q(\STAGEN[38].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[311]),
        .Q(\STAGEN[38].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__36_n_0),
        .Q(\STAGEN[38].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__36_n_0),
        .Q(\STAGEN[38].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__36_n_0),
        .Q(w_bit_up_39),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_38),
        .Q(\STAGEN[38].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[38].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_39),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__36_n_0),
        .Q(\STAGEN[38].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_38),
        .Q(\STAGEN[38].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[38].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[38].stage/split_module/p_1_out ),
        .Q(w_swap_up_39),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[0]_i_1__38_n_0 ),
        .Q(readdata_o[312]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[1]_i_1__38_n_0 ),
        .Q(readdata_o[313]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[2]_i_1__38_n_0 ),
        .Q(readdata_o[314]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[3]_i_1__38_n_0 ),
        .Q(readdata_o[315]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[4]_i_1__38_n_0 ),
        .Q(readdata_o[316]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[5]_i_1__38_n_0 ),
        .Q(readdata_o[317]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[6]_i_1__38_n_0 ),
        .Q(readdata_o[318]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__38_n_0 ),
        .D(\r_data[7]_i_2__38_n_0 ),
        .Q(readdata_o[319]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_39),
        .Q(\STAGEN[39].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[319]),
        .Q(\STAGEN[39].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__37_n_0),
        .Q(\STAGEN[39].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__37_n_0),
        .Q(\STAGEN[39].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__37_n_0),
        .Q(w_bit_up_40),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_39),
        .Q(\STAGEN[39].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[39].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_40),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__37_n_0),
        .Q(\STAGEN[39].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_39),
        .Q(\STAGEN[39].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[39].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[39].stage/split_module/p_1_out ),
        .Q(w_swap_up_40),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[0]_i_1__2_n_0 ),
        .Q(readdata_o[24]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[1]_i_1__2_n_0 ),
        .Q(readdata_o[25]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[2]_i_1__2_n_0 ),
        .Q(readdata_o[26]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[3]_i_1__2_n_0 ),
        .Q(readdata_o[27]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[4]_i_1__2_n_0 ),
        .Q(readdata_o[28]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[5]_i_1__2_n_0 ),
        .Q(readdata_o[29]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[6]_i_1__2_n_0 ),
        .Q(readdata_o[30]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__2_n_0 ),
        .D(\r_data[7]_i_2__2_n_0 ),
        .Q(readdata_o[31]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_3),
        .Q(\STAGEN[3].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[31]),
        .Q(\STAGEN[3].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__1_n_0),
        .Q(\STAGEN[3].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__1_n_0),
        .Q(\STAGEN[3].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__1_n_0),
        .Q(w_bit_up_4),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_3),
        .Q(\STAGEN[3].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[3].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_4),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__1_n_0),
        .Q(\STAGEN[3].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_3),
        .Q(\STAGEN[3].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[3].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[3].stage/split_module/p_1_out ),
        .Q(w_swap_up_4),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[0]_i_1__39_n_0 ),
        .Q(readdata_o[320]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[1]_i_1__39_n_0 ),
        .Q(readdata_o[321]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[2]_i_1__39_n_0 ),
        .Q(readdata_o[322]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[3]_i_1__39_n_0 ),
        .Q(readdata_o[323]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[4]_i_1__39_n_0 ),
        .Q(readdata_o[324]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[5]_i_1__39_n_0 ),
        .Q(readdata_o[325]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[6]_i_1__39_n_0 ),
        .Q(readdata_o[326]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__39_n_0 ),
        .D(\r_data[7]_i_2__39_n_0 ),
        .Q(readdata_o[327]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_40),
        .Q(\STAGEN[40].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[327]),
        .Q(\STAGEN[40].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__38_n_0),
        .Q(\STAGEN[40].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__38_n_0),
        .Q(\STAGEN[40].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__38_n_0),
        .Q(w_bit_up_41),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_40),
        .Q(\STAGEN[40].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[40].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_41),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__38_n_0),
        .Q(\STAGEN[40].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_40),
        .Q(\STAGEN[40].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[40].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[40].stage/split_module/p_1_out ),
        .Q(w_swap_up_41),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[0]_i_1__40_n_0 ),
        .Q(readdata_o[328]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[1]_i_1__40_n_0 ),
        .Q(readdata_o[329]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[2]_i_1__40_n_0 ),
        .Q(readdata_o[330]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[3]_i_1__40_n_0 ),
        .Q(readdata_o[331]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[4]_i_1__40_n_0 ),
        .Q(readdata_o[332]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[5]_i_1__40_n_0 ),
        .Q(readdata_o[333]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[6]_i_1__40_n_0 ),
        .Q(readdata_o[334]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__40_n_0 ),
        .D(\r_data[7]_i_2__40_n_0 ),
        .Q(readdata_o[335]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_41),
        .Q(\STAGEN[41].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[335]),
        .Q(\STAGEN[41].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__39_n_0),
        .Q(\STAGEN[41].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__39_n_0),
        .Q(\STAGEN[41].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__39_n_0),
        .Q(w_bit_up_42),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_41),
        .Q(\STAGEN[41].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[41].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_42),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__39_n_0),
        .Q(\STAGEN[41].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_41),
        .Q(\STAGEN[41].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[41].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[41].stage/split_module/p_1_out ),
        .Q(w_swap_up_42),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[0]_i_1__41_n_0 ),
        .Q(readdata_o[336]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[1]_i_1__41_n_0 ),
        .Q(readdata_o[337]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[2]_i_1__41_n_0 ),
        .Q(readdata_o[338]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[3]_i_1__41_n_0 ),
        .Q(readdata_o[339]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[4]_i_1__41_n_0 ),
        .Q(readdata_o[340]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[5]_i_1__41_n_0 ),
        .Q(readdata_o[341]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[6]_i_1__41_n_0 ),
        .Q(readdata_o[342]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__41_n_0 ),
        .D(\r_data[7]_i_2__41_n_0 ),
        .Q(readdata_o[343]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_42),
        .Q(\STAGEN[42].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[343]),
        .Q(\STAGEN[42].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__40_n_0),
        .Q(\STAGEN[42].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__40_n_0),
        .Q(\STAGEN[42].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__40_n_0),
        .Q(w_bit_up_43),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_42),
        .Q(\STAGEN[42].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[42].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_43),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__40_n_0),
        .Q(\STAGEN[42].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_42),
        .Q(\STAGEN[42].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[42].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[42].stage/split_module/p_1_out ),
        .Q(w_swap_up_43),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[0]_i_1__42_n_0 ),
        .Q(readdata_o[344]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[1]_i_1__42_n_0 ),
        .Q(readdata_o[345]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[2]_i_1__42_n_0 ),
        .Q(readdata_o[346]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[3]_i_1__42_n_0 ),
        .Q(readdata_o[347]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[4]_i_1__42_n_0 ),
        .Q(readdata_o[348]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[5]_i_1__42_n_0 ),
        .Q(readdata_o[349]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[6]_i_1__42_n_0 ),
        .Q(readdata_o[350]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__42_n_0 ),
        .D(\r_data[7]_i_2__42_n_0 ),
        .Q(readdata_o[351]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_43),
        .Q(\STAGEN[43].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[351]),
        .Q(\STAGEN[43].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__41_n_0),
        .Q(\STAGEN[43].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__41_n_0),
        .Q(\STAGEN[43].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__41_n_0),
        .Q(w_bit_up_44),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_43),
        .Q(\STAGEN[43].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[43].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_44),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__41_n_0),
        .Q(\STAGEN[43].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_43),
        .Q(\STAGEN[43].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[43].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[43].stage/split_module/p_1_out ),
        .Q(w_swap_up_44),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[0]_i_1__43_n_0 ),
        .Q(readdata_o[352]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[1]_i_1__43_n_0 ),
        .Q(readdata_o[353]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[2]_i_1__43_n_0 ),
        .Q(readdata_o[354]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[3]_i_1__43_n_0 ),
        .Q(readdata_o[355]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[4]_i_1__43_n_0 ),
        .Q(readdata_o[356]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[5]_i_1__43_n_0 ),
        .Q(readdata_o[357]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[6]_i_1__43_n_0 ),
        .Q(readdata_o[358]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__43_n_0 ),
        .D(\r_data[7]_i_2__43_n_0 ),
        .Q(readdata_o[359]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_44),
        .Q(\STAGEN[44].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[359]),
        .Q(\STAGEN[44].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__42_n_0),
        .Q(\STAGEN[44].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__42_n_0),
        .Q(\STAGEN[44].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__42_n_0),
        .Q(w_bit_up_45),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_44),
        .Q(\STAGEN[44].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[44].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_45),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__42_n_0),
        .Q(\STAGEN[44].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_44),
        .Q(\STAGEN[44].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[44].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[44].stage/split_module/p_1_out ),
        .Q(w_swap_up_45),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[0]_i_1__44_n_0 ),
        .Q(readdata_o[360]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[1]_i_1__44_n_0 ),
        .Q(readdata_o[361]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[2]_i_1__44_n_0 ),
        .Q(readdata_o[362]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[3]_i_1__44_n_0 ),
        .Q(readdata_o[363]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[4]_i_1__44_n_0 ),
        .Q(readdata_o[364]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[5]_i_1__44_n_0 ),
        .Q(readdata_o[365]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[6]_i_1__44_n_0 ),
        .Q(readdata_o[366]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__44_n_0 ),
        .D(\r_data[7]_i_2__44_n_0 ),
        .Q(readdata_o[367]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_45),
        .Q(\STAGEN[45].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[367]),
        .Q(\STAGEN[45].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__43_n_0),
        .Q(\STAGEN[45].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__43_n_0),
        .Q(\STAGEN[45].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__43_n_0),
        .Q(w_bit_up_46),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_45),
        .Q(\STAGEN[45].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[45].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_46),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__43_n_0),
        .Q(\STAGEN[45].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_45),
        .Q(\STAGEN[45].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[45].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[45].stage/split_module/p_1_out ),
        .Q(w_swap_up_46),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[0]_i_1__45_n_0 ),
        .Q(readdata_o[368]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[1]_i_1__45_n_0 ),
        .Q(readdata_o[369]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[2]_i_1__45_n_0 ),
        .Q(readdata_o[370]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[3]_i_1__45_n_0 ),
        .Q(readdata_o[371]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[4]_i_1__45_n_0 ),
        .Q(readdata_o[372]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[5]_i_1__45_n_0 ),
        .Q(readdata_o[373]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[6]_i_1__45_n_0 ),
        .Q(readdata_o[374]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__45_n_0 ),
        .D(\r_data[7]_i_2__45_n_0 ),
        .Q(readdata_o[375]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_46),
        .Q(\STAGEN[46].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[375]),
        .Q(\STAGEN[46].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__44_n_0),
        .Q(\STAGEN[46].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__44_n_0),
        .Q(\STAGEN[46].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__44_n_0),
        .Q(w_bit_up_47),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_46),
        .Q(\STAGEN[46].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[46].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_47),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__44_n_0),
        .Q(\STAGEN[46].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_46),
        .Q(\STAGEN[46].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[46].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[46].stage/split_module/p_1_out ),
        .Q(w_swap_up_47),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[0]_i_1__46_n_0 ),
        .Q(readdata_o[376]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[1]_i_1__46_n_0 ),
        .Q(readdata_o[377]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[2]_i_1__46_n_0 ),
        .Q(readdata_o[378]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[3]_i_1__46_n_0 ),
        .Q(readdata_o[379]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[4]_i_1__46_n_0 ),
        .Q(readdata_o[380]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[5]_i_1__46_n_0 ),
        .Q(readdata_o[381]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[6]_i_1__46_n_0 ),
        .Q(readdata_o[382]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__46_n_0 ),
        .D(\r_data[7]_i_2__46_n_0 ),
        .Q(readdata_o[383]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_47),
        .Q(\STAGEN[47].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[383]),
        .Q(\STAGEN[47].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__45_n_0),
        .Q(\STAGEN[47].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__45_n_0),
        .Q(\STAGEN[47].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__45_n_0),
        .Q(w_bit_up_48),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_47),
        .Q(\STAGEN[47].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[47].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_48),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__45_n_0),
        .Q(\STAGEN[47].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_47),
        .Q(\STAGEN[47].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[47].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[47].stage/split_module/p_1_out ),
        .Q(w_swap_up_48),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[0]_i_1__47_n_0 ),
        .Q(readdata_o[384]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[1]_i_1__47_n_0 ),
        .Q(readdata_o[385]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[2]_i_1__47_n_0 ),
        .Q(readdata_o[386]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[3]_i_1__47_n_0 ),
        .Q(readdata_o[387]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[4]_i_1__47_n_0 ),
        .Q(readdata_o[388]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[5]_i_1__47_n_0 ),
        .Q(readdata_o[389]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[6]_i_1__47_n_0 ),
        .Q(readdata_o[390]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__47_n_0 ),
        .D(\r_data[7]_i_2__47_n_0 ),
        .Q(readdata_o[391]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_48),
        .Q(\STAGEN[48].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[391]),
        .Q(\STAGEN[48].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__46_n_0),
        .Q(\STAGEN[48].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__46_n_0),
        .Q(\STAGEN[48].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_48),
        .Q(\STAGEN[48].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[48].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_49),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__46_n_0),
        .Q(\STAGEN[48].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_48),
        .Q(\STAGEN[48].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[48].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[48].stage/split_module/p_1_out ),
        .Q(\STAGEN[48].stage/split_module/r_swap_reg_n_0_[1] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[0]_i_1__3_n_0 ),
        .Q(readdata_o[32]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[1]_i_1__3_n_0 ),
        .Q(readdata_o[33]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[2]_i_1__3_n_0 ),
        .Q(readdata_o[34]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[3]_i_1__3_n_0 ),
        .Q(readdata_o[35]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[4]_i_1__3_n_0 ),
        .Q(readdata_o[36]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[5]_i_1__3_n_0 ),
        .Q(readdata_o[37]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[6]_i_1__3_n_0 ),
        .Q(readdata_o[38]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__3_n_0 ),
        .D(\r_data[7]_i_2__3_n_0 ),
        .Q(readdata_o[39]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_4),
        .Q(\STAGEN[4].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[39]),
        .Q(\STAGEN[4].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__2_n_0),
        .Q(\STAGEN[4].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__2_n_0),
        .Q(\STAGEN[4].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__2_n_0),
        .Q(w_bit_up_5),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_4),
        .Q(\STAGEN[4].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[4].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_5),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__2_n_0),
        .Q(\STAGEN[4].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_4),
        .Q(\STAGEN[4].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[4].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[4].stage/split_module/p_1_out ),
        .Q(w_swap_up_5),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[0]_i_1__4_n_0 ),
        .Q(readdata_o[40]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[1]_i_1__4_n_0 ),
        .Q(readdata_o[41]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[2]_i_1__4_n_0 ),
        .Q(readdata_o[42]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[3]_i_1__4_n_0 ),
        .Q(readdata_o[43]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[4]_i_1__4_n_0 ),
        .Q(readdata_o[44]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[5]_i_1__4_n_0 ),
        .Q(readdata_o[45]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[6]_i_1__4_n_0 ),
        .Q(readdata_o[46]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__4_n_0 ),
        .D(\r_data[7]_i_2__4_n_0 ),
        .Q(readdata_o[47]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_5),
        .Q(\STAGEN[5].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[47]),
        .Q(\STAGEN[5].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__3_n_0),
        .Q(\STAGEN[5].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__3_n_0),
        .Q(\STAGEN[5].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__3_n_0),
        .Q(w_bit_up_6),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_5),
        .Q(\STAGEN[5].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[5].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_6),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__3_n_0),
        .Q(\STAGEN[5].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_5),
        .Q(\STAGEN[5].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[5].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[5].stage/split_module/p_1_out ),
        .Q(w_swap_up_6),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[0]_i_1__5_n_0 ),
        .Q(readdata_o[48]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[1]_i_1__5_n_0 ),
        .Q(readdata_o[49]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[2]_i_1__5_n_0 ),
        .Q(readdata_o[50]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[3]_i_1__5_n_0 ),
        .Q(readdata_o[51]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[4]_i_1__5_n_0 ),
        .Q(readdata_o[52]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[5]_i_1__5_n_0 ),
        .Q(readdata_o[53]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[6]_i_1__5_n_0 ),
        .Q(readdata_o[54]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__5_n_0 ),
        .D(\r_data[7]_i_2__5_n_0 ),
        .Q(readdata_o[55]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_6),
        .Q(\STAGEN[6].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[55]),
        .Q(\STAGEN[6].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__4_n_0),
        .Q(\STAGEN[6].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__4_n_0),
        .Q(\STAGEN[6].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__4_n_0),
        .Q(w_bit_up_7),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_6),
        .Q(\STAGEN[6].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[6].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_7),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__4_n_0),
        .Q(\STAGEN[6].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_6),
        .Q(\STAGEN[6].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[6].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[6].stage/split_module/p_1_out ),
        .Q(w_swap_up_7),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[0]_i_1__6_n_0 ),
        .Q(readdata_o[56]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[1]_i_1__6_n_0 ),
        .Q(readdata_o[57]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[2]_i_1__6_n_0 ),
        .Q(readdata_o[58]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[3]_i_1__6_n_0 ),
        .Q(readdata_o[59]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[4]_i_1__6_n_0 ),
        .Q(readdata_o[60]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[5]_i_1__6_n_0 ),
        .Q(readdata_o[61]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[6]_i_1__6_n_0 ),
        .Q(readdata_o[62]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__6_n_0 ),
        .D(\r_data[7]_i_2__6_n_0 ),
        .Q(readdata_o[63]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_7),
        .Q(\STAGEN[7].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[63]),
        .Q(\STAGEN[7].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__5_n_0),
        .Q(\STAGEN[7].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__5_n_0),
        .Q(\STAGEN[7].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__5_n_0),
        .Q(w_bit_up_8),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_7),
        .Q(\STAGEN[7].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[7].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_8),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__5_n_0),
        .Q(\STAGEN[7].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_7),
        .Q(\STAGEN[7].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[7].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[7].stage/split_module/p_1_out ),
        .Q(w_swap_up_8),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[0]_i_1__7_n_0 ),
        .Q(readdata_o[64]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[1]_i_1__7_n_0 ),
        .Q(readdata_o[65]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[2]_i_1__7_n_0 ),
        .Q(readdata_o[66]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[3]_i_1__7_n_0 ),
        .Q(readdata_o[67]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[4]_i_1__7_n_0 ),
        .Q(readdata_o[68]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[5]_i_1__7_n_0 ),
        .Q(readdata_o[69]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[6]_i_1__7_n_0 ),
        .Q(readdata_o[70]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__7_n_0 ),
        .D(\r_data[7]_i_2__7_n_0 ),
        .Q(readdata_o[71]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_8),
        .Q(\STAGEN[8].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[71]),
        .Q(\STAGEN[8].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__6_n_0),
        .Q(\STAGEN[8].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__6_n_0),
        .Q(\STAGEN[8].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__6_n_0),
        .Q(w_bit_up_9),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_8),
        .Q(\STAGEN[8].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[8].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_9),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__6_n_0),
        .Q(\STAGEN[8].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_8),
        .Q(\STAGEN[8].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[8].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[8].stage/split_module/p_1_out ),
        .Q(w_swap_up_9),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[0] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[0]_i_1__8_n_0 ),
        .Q(readdata_o[72]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[1] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[1]_i_1__8_n_0 ),
        .Q(readdata_o[73]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[2] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[2]_i_1__8_n_0 ),
        .Q(readdata_o[74]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[3] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[3]_i_1__8_n_0 ),
        .Q(readdata_o[75]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[4] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[4]_i_1__8_n_0 ),
        .Q(readdata_o[76]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[5] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[5]_i_1__8_n_0 ),
        .Q(readdata_o[77]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[6] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[6]_i_1__8_n_0 ),
        .Q(readdata_o[78]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/r_data_reg[7] 
       (.C(clk),
        .CE(\r_data[7]_i_1__8_n_0 ),
        .D(\r_data[7]_i_2__8_n_0 ),
        .Q(readdata_o[79]),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_bit1_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_bit_up_9),
        .Q(\STAGEN[9].stage/split_module/r_bit1 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_bit2_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(readdata_o[79]),
        .Q(\STAGEN[9].stage/split_module/r_bit2 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_compare_result_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_compare_result_i_1__7_n_0),
        .Q(\STAGEN[9].stage/split_module/r_compare_result ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_freeze_compare_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_freeze_compare_i_1__7_n_0),
        .Q(\STAGEN[9].stage/split_module/r_freeze_compare_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_large_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_large_bit_i_1__7_n_0),
        .Q(w_bit_up_10),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_run_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_9),
        .Q(\STAGEN[9].stage/split_module/r_run_reg_n_0_[0] ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_run_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[9].stage/split_module/r_run_reg_n_0_[0] ),
        .Q(w_run_up_10),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_small_bit_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_small_bit_i_1__7_n_0),
        .Q(\STAGEN[9].stage/split_module/r_small_bit_reg_n_0 ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_swap_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_swap_up_9),
        .Q(\STAGEN[9].stage/split_module/p_0_in ),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \STAGEN[9].stage/split_module/r_swap_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[9].stage/split_module/p_1_out ),
        .Q(w_swap_up_10),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  VCC VCC
       (.P(\<const1>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_done_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_done_i_1_n_0),
        .Q(done_o),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[0] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(r_pulses0),
        .Q(\interrupt_module/r_pulses_reg_n_0_ ),
        .S(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[1] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(r_pulses),
        .Q(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .R(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[2] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(\r_pulses[2]_i_1_n_0 ),
        .Q(\interrupt_module/r_pulses_reg_n_0_[2] ),
        .R(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDSE #(
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_S_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[3] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(\r_pulses[3]_i_1_n_0 ),
        .Q(\interrupt_module/r_pulses_reg_n_0_[3] ),
        .S(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[4] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(\r_pulses[4]_i_1_n_0 ),
        .Q(\interrupt_module/r_pulses_reg_n_0_[4] ),
        .R(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_pulses_reg[5] 
       (.C(clk),
        .CE(\r_pulses[5]_i_2_n_0 ),
        .D(\r_pulses[5]_i_3_n_0 ),
        .Q(interrupt_o),
        .R(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_run_delay_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_49),
        .Q(\interrupt_module/r_run_delay ),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \interrupt_module/r_swap_delay_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\STAGEN[48].stage/split_module/r_swap_reg_n_0_[1] ),
        .Q(\interrupt_module/r_swap_delay ),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1
       (.I0(readdata_o[15]),
        .I1(w_bit_up_1),
        .I2(\STAGEN[1].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[1].stage/split_module/r_compare_result ),
        .I4(w_run_up_1),
        .O(r_compare_result_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__0
       (.I0(readdata_o[23]),
        .I1(w_bit_up_2),
        .I2(\STAGEN[2].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[2].stage/split_module/r_compare_result ),
        .I4(w_run_up_2),
        .O(r_compare_result_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__1
       (.I0(readdata_o[31]),
        .I1(w_bit_up_3),
        .I2(\STAGEN[3].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[3].stage/split_module/r_compare_result ),
        .I4(w_run_up_3),
        .O(r_compare_result_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__10
       (.I0(readdata_o[103]),
        .I1(w_bit_up_12),
        .I2(\STAGEN[12].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[12].stage/split_module/r_compare_result ),
        .I4(w_run_up_12),
        .O(r_compare_result_i_1__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__11
       (.I0(readdata_o[111]),
        .I1(w_bit_up_13),
        .I2(\STAGEN[13].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[13].stage/split_module/r_compare_result ),
        .I4(w_run_up_13),
        .O(r_compare_result_i_1__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__12
       (.I0(readdata_o[119]),
        .I1(w_bit_up_14),
        .I2(\STAGEN[14].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[14].stage/split_module/r_compare_result ),
        .I4(w_run_up_14),
        .O(r_compare_result_i_1__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__13
       (.I0(readdata_o[127]),
        .I1(w_bit_up_15),
        .I2(\STAGEN[15].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[15].stage/split_module/r_compare_result ),
        .I4(w_run_up_15),
        .O(r_compare_result_i_1__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__14
       (.I0(readdata_o[135]),
        .I1(w_bit_up_16),
        .I2(\STAGEN[16].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[16].stage/split_module/r_compare_result ),
        .I4(w_run_up_16),
        .O(r_compare_result_i_1__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__15
       (.I0(readdata_o[143]),
        .I1(w_bit_up_17),
        .I2(\STAGEN[17].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[17].stage/split_module/r_compare_result ),
        .I4(w_run_up_17),
        .O(r_compare_result_i_1__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__16
       (.I0(readdata_o[151]),
        .I1(w_bit_up_18),
        .I2(\STAGEN[18].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[18].stage/split_module/r_compare_result ),
        .I4(w_run_up_18),
        .O(r_compare_result_i_1__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__17
       (.I0(readdata_o[159]),
        .I1(w_bit_up_19),
        .I2(\STAGEN[19].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[19].stage/split_module/r_compare_result ),
        .I4(w_run_up_19),
        .O(r_compare_result_i_1__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__18
       (.I0(readdata_o[167]),
        .I1(w_bit_up_20),
        .I2(\STAGEN[20].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[20].stage/split_module/r_compare_result ),
        .I4(w_run_up_20),
        .O(r_compare_result_i_1__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__19
       (.I0(readdata_o[175]),
        .I1(w_bit_up_21),
        .I2(\STAGEN[21].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[21].stage/split_module/r_compare_result ),
        .I4(w_run_up_21),
        .O(r_compare_result_i_1__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__2
       (.I0(readdata_o[39]),
        .I1(w_bit_up_4),
        .I2(\STAGEN[4].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[4].stage/split_module/r_compare_result ),
        .I4(w_run_up_4),
        .O(r_compare_result_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__20
       (.I0(readdata_o[183]),
        .I1(w_bit_up_22),
        .I2(\STAGEN[22].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[22].stage/split_module/r_compare_result ),
        .I4(w_run_up_22),
        .O(r_compare_result_i_1__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__21
       (.I0(readdata_o[191]),
        .I1(w_bit_up_23),
        .I2(\STAGEN[23].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[23].stage/split_module/r_compare_result ),
        .I4(w_run_up_23),
        .O(r_compare_result_i_1__21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__22
       (.I0(readdata_o[199]),
        .I1(w_bit_up_24),
        .I2(\STAGEN[24].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[24].stage/split_module/r_compare_result ),
        .I4(w_run_up_24),
        .O(r_compare_result_i_1__22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__23
       (.I0(readdata_o[207]),
        .I1(w_bit_up_25),
        .I2(\STAGEN[25].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[25].stage/split_module/r_compare_result ),
        .I4(w_run_up_25),
        .O(r_compare_result_i_1__23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__24
       (.I0(readdata_o[215]),
        .I1(w_bit_up_26),
        .I2(\STAGEN[26].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[26].stage/split_module/r_compare_result ),
        .I4(w_run_up_26),
        .O(r_compare_result_i_1__24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__25
       (.I0(readdata_o[223]),
        .I1(w_bit_up_27),
        .I2(\STAGEN[27].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[27].stage/split_module/r_compare_result ),
        .I4(w_run_up_27),
        .O(r_compare_result_i_1__25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__26
       (.I0(readdata_o[231]),
        .I1(w_bit_up_28),
        .I2(\STAGEN[28].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[28].stage/split_module/r_compare_result ),
        .I4(w_run_up_28),
        .O(r_compare_result_i_1__26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__27
       (.I0(readdata_o[239]),
        .I1(w_bit_up_29),
        .I2(\STAGEN[29].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[29].stage/split_module/r_compare_result ),
        .I4(w_run_up_29),
        .O(r_compare_result_i_1__27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__28
       (.I0(readdata_o[247]),
        .I1(w_bit_up_30),
        .I2(\STAGEN[30].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[30].stage/split_module/r_compare_result ),
        .I4(w_run_up_30),
        .O(r_compare_result_i_1__28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__29
       (.I0(readdata_o[255]),
        .I1(w_bit_up_31),
        .I2(\STAGEN[31].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[31].stage/split_module/r_compare_result ),
        .I4(w_run_up_31),
        .O(r_compare_result_i_1__29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__3
       (.I0(readdata_o[47]),
        .I1(w_bit_up_5),
        .I2(\STAGEN[5].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[5].stage/split_module/r_compare_result ),
        .I4(w_run_up_5),
        .O(r_compare_result_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__30
       (.I0(readdata_o[263]),
        .I1(w_bit_up_32),
        .I2(\STAGEN[32].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[32].stage/split_module/r_compare_result ),
        .I4(w_run_up_32),
        .O(r_compare_result_i_1__30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__31
       (.I0(readdata_o[271]),
        .I1(w_bit_up_33),
        .I2(\STAGEN[33].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[33].stage/split_module/r_compare_result ),
        .I4(w_run_up_33),
        .O(r_compare_result_i_1__31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__32
       (.I0(readdata_o[279]),
        .I1(w_bit_up_34),
        .I2(\STAGEN[34].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[34].stage/split_module/r_compare_result ),
        .I4(w_run_up_34),
        .O(r_compare_result_i_1__32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__33
       (.I0(readdata_o[287]),
        .I1(w_bit_up_35),
        .I2(\STAGEN[35].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[35].stage/split_module/r_compare_result ),
        .I4(w_run_up_35),
        .O(r_compare_result_i_1__33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__34
       (.I0(readdata_o[295]),
        .I1(w_bit_up_36),
        .I2(\STAGEN[36].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[36].stage/split_module/r_compare_result ),
        .I4(w_run_up_36),
        .O(r_compare_result_i_1__34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__35
       (.I0(readdata_o[303]),
        .I1(w_bit_up_37),
        .I2(\STAGEN[37].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[37].stage/split_module/r_compare_result ),
        .I4(w_run_up_37),
        .O(r_compare_result_i_1__35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__36
       (.I0(readdata_o[311]),
        .I1(w_bit_up_38),
        .I2(\STAGEN[38].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[38].stage/split_module/r_compare_result ),
        .I4(w_run_up_38),
        .O(r_compare_result_i_1__36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__37
       (.I0(readdata_o[319]),
        .I1(w_bit_up_39),
        .I2(\STAGEN[39].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[39].stage/split_module/r_compare_result ),
        .I4(w_run_up_39),
        .O(r_compare_result_i_1__37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__38
       (.I0(readdata_o[327]),
        .I1(w_bit_up_40),
        .I2(\STAGEN[40].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[40].stage/split_module/r_compare_result ),
        .I4(w_run_up_40),
        .O(r_compare_result_i_1__38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__39
       (.I0(readdata_o[335]),
        .I1(w_bit_up_41),
        .I2(\STAGEN[41].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[41].stage/split_module/r_compare_result ),
        .I4(w_run_up_41),
        .O(r_compare_result_i_1__39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__4
       (.I0(readdata_o[55]),
        .I1(w_bit_up_6),
        .I2(\STAGEN[6].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[6].stage/split_module/r_compare_result ),
        .I4(w_run_up_6),
        .O(r_compare_result_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__40
       (.I0(readdata_o[343]),
        .I1(w_bit_up_42),
        .I2(\STAGEN[42].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[42].stage/split_module/r_compare_result ),
        .I4(w_run_up_42),
        .O(r_compare_result_i_1__40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__41
       (.I0(readdata_o[351]),
        .I1(w_bit_up_43),
        .I2(\STAGEN[43].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[43].stage/split_module/r_compare_result ),
        .I4(w_run_up_43),
        .O(r_compare_result_i_1__41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__42
       (.I0(readdata_o[359]),
        .I1(w_bit_up_44),
        .I2(\STAGEN[44].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[44].stage/split_module/r_compare_result ),
        .I4(w_run_up_44),
        .O(r_compare_result_i_1__42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__43
       (.I0(readdata_o[367]),
        .I1(w_bit_up_45),
        .I2(\STAGEN[45].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[45].stage/split_module/r_compare_result ),
        .I4(w_run_up_45),
        .O(r_compare_result_i_1__43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__44
       (.I0(readdata_o[375]),
        .I1(w_bit_up_46),
        .I2(\STAGEN[46].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[46].stage/split_module/r_compare_result ),
        .I4(w_run_up_46),
        .O(r_compare_result_i_1__44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__45
       (.I0(readdata_o[383]),
        .I1(w_bit_up_47),
        .I2(\STAGEN[47].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[47].stage/split_module/r_compare_result ),
        .I4(w_run_up_47),
        .O(r_compare_result_i_1__45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__46
       (.I0(readdata_o[391]),
        .I1(w_bit_up_48),
        .I2(\STAGEN[48].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[48].stage/split_module/r_compare_result ),
        .I4(w_run_up_48),
        .O(r_compare_result_i_1__46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__5
       (.I0(readdata_o[63]),
        .I1(w_bit_up_7),
        .I2(\STAGEN[7].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[7].stage/split_module/r_compare_result ),
        .I4(w_run_up_7),
        .O(r_compare_result_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__6
       (.I0(readdata_o[71]),
        .I1(w_bit_up_8),
        .I2(\STAGEN[8].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[8].stage/split_module/r_compare_result ),
        .I4(w_run_up_8),
        .O(r_compare_result_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__7
       (.I0(readdata_o[79]),
        .I1(w_bit_up_9),
        .I2(\STAGEN[9].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[9].stage/split_module/r_compare_result ),
        .I4(w_run_up_9),
        .O(r_compare_result_i_1__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__8
       (.I0(readdata_o[87]),
        .I1(w_bit_up_10),
        .I2(\STAGEN[10].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[10].stage/split_module/r_compare_result ),
        .I4(w_run_up_10),
        .O(r_compare_result_i_1__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT5 #(
    .INIT(32'hF4040000)) 
    r_compare_result_i_1__9
       (.I0(readdata_o[95]),
        .I1(w_bit_up_11),
        .I2(\STAGEN[11].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I3(\STAGEN[11].stage/split_module/r_compare_result ),
        .I4(w_run_up_11),
        .O(r_compare_result_i_1__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_count[3]_i_1 
       (.I0(start_i),
        .I1(rst),
        .O(r_count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1 
       (.I0(writedata_i[0]),
        .I1(r_small_bit),
        .I2(load_i[0]),
        .O(\r_data[0]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__0 
       (.I0(writedata_i[8]),
        .I1(\STAGEN[2].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[1]),
        .O(r_data));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__1 
       (.I0(writedata_i[16]),
        .I1(\STAGEN[3].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[2]),
        .O(\r_data[0]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__10 
       (.I0(writedata_i[88]),
        .I1(\STAGEN[12].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[11]),
        .O(\r_data[0]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__11 
       (.I0(writedata_i[96]),
        .I1(\STAGEN[13].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[12]),
        .O(\r_data[0]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__12 
       (.I0(writedata_i[104]),
        .I1(\STAGEN[14].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[13]),
        .O(\r_data[0]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__13 
       (.I0(writedata_i[112]),
        .I1(\STAGEN[15].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[14]),
        .O(\r_data[0]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__14 
       (.I0(writedata_i[120]),
        .I1(\STAGEN[16].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[15]),
        .O(\r_data[0]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__15 
       (.I0(writedata_i[128]),
        .I1(\STAGEN[17].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[16]),
        .O(\r_data[0]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__16 
       (.I0(writedata_i[136]),
        .I1(\STAGEN[18].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[17]),
        .O(\r_data[0]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__17 
       (.I0(writedata_i[144]),
        .I1(\STAGEN[19].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[18]),
        .O(\r_data[0]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__18 
       (.I0(writedata_i[152]),
        .I1(\STAGEN[20].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[19]),
        .O(\r_data[0]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__19 
       (.I0(writedata_i[160]),
        .I1(\STAGEN[21].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[20]),
        .O(\r_data[0]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__2 
       (.I0(writedata_i[24]),
        .I1(\STAGEN[4].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[3]),
        .O(\r_data[0]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__20 
       (.I0(writedata_i[168]),
        .I1(\STAGEN[22].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[21]),
        .O(\r_data[0]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__21 
       (.I0(writedata_i[176]),
        .I1(\STAGEN[23].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[22]),
        .O(\r_data[0]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__22 
       (.I0(writedata_i[184]),
        .I1(\STAGEN[24].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[23]),
        .O(\r_data[0]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__23 
       (.I0(writedata_i[192]),
        .I1(\STAGEN[25].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[24]),
        .O(\r_data[0]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__24 
       (.I0(writedata_i[200]),
        .I1(\STAGEN[26].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[25]),
        .O(\r_data[0]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__25 
       (.I0(writedata_i[208]),
        .I1(\STAGEN[27].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[26]),
        .O(\r_data[0]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__26 
       (.I0(writedata_i[216]),
        .I1(\STAGEN[28].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[27]),
        .O(\r_data[0]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__27 
       (.I0(writedata_i[224]),
        .I1(\STAGEN[29].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[28]),
        .O(\r_data[0]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__28 
       (.I0(writedata_i[232]),
        .I1(\STAGEN[30].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[29]),
        .O(\r_data[0]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__29 
       (.I0(writedata_i[240]),
        .I1(\STAGEN[31].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[30]),
        .O(\r_data[0]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__3 
       (.I0(writedata_i[32]),
        .I1(\STAGEN[5].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[4]),
        .O(\r_data[0]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__30 
       (.I0(writedata_i[248]),
        .I1(\STAGEN[32].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[31]),
        .O(\r_data[0]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__31 
       (.I0(writedata_i[256]),
        .I1(\STAGEN[33].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[32]),
        .O(\r_data[0]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__32 
       (.I0(writedata_i[264]),
        .I1(\STAGEN[34].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[33]),
        .O(\r_data[0]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__33 
       (.I0(writedata_i[272]),
        .I1(\STAGEN[35].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[34]),
        .O(\r_data[0]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__34 
       (.I0(writedata_i[280]),
        .I1(\STAGEN[36].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[35]),
        .O(\r_data[0]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__35 
       (.I0(writedata_i[288]),
        .I1(\STAGEN[37].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[36]),
        .O(\r_data[0]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__36 
       (.I0(writedata_i[296]),
        .I1(\STAGEN[38].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[37]),
        .O(\r_data[0]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__37 
       (.I0(writedata_i[304]),
        .I1(\STAGEN[39].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[38]),
        .O(\r_data[0]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__38 
       (.I0(writedata_i[312]),
        .I1(\STAGEN[40].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[39]),
        .O(\r_data[0]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__39 
       (.I0(writedata_i[320]),
        .I1(\STAGEN[41].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[40]),
        .O(\r_data[0]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__4 
       (.I0(writedata_i[40]),
        .I1(\STAGEN[6].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[5]),
        .O(\r_data[0]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__40 
       (.I0(writedata_i[328]),
        .I1(\STAGEN[42].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[41]),
        .O(\r_data[0]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__41 
       (.I0(writedata_i[336]),
        .I1(\STAGEN[43].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[42]),
        .O(\r_data[0]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__42 
       (.I0(writedata_i[344]),
        .I1(\STAGEN[44].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[43]),
        .O(\r_data[0]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__43 
       (.I0(writedata_i[352]),
        .I1(\STAGEN[45].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[44]),
        .O(\r_data[0]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__44 
       (.I0(writedata_i[360]),
        .I1(\STAGEN[46].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[45]),
        .O(\r_data[0]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__45 
       (.I0(writedata_i[368]),
        .I1(\STAGEN[47].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[46]),
        .O(\r_data[0]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__46 
       (.I0(writedata_i[376]),
        .I1(\STAGEN[48].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[47]),
        .O(\r_data[0]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__47 
       (.I0(writedata_i[384]),
        .I1(r_value_66),
        .I2(load_i[48]),
        .O(\r_data[0]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__5 
       (.I0(writedata_i[48]),
        .I1(\STAGEN[7].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[6]),
        .O(\r_data[0]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__6 
       (.I0(writedata_i[56]),
        .I1(\STAGEN[8].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[7]),
        .O(\r_data[0]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__7 
       (.I0(writedata_i[64]),
        .I1(\STAGEN[9].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[8]),
        .O(\r_data[0]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__8 
       (.I0(writedata_i[72]),
        .I1(\STAGEN[10].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[9]),
        .O(\r_data[0]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[0]_i_1__9 
       (.I0(writedata_i[80]),
        .I1(\STAGEN[11].stage/split_module/r_small_bit_reg_n_0 ),
        .I2(load_i[10]),
        .O(\r_data[0]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1 
       (.I0(writedata_i[1]),
        .I1(readdata_o[0]),
        .I2(load_i[0]),
        .O(\r_data[1]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__0 
       (.I0(writedata_i[9]),
        .I1(readdata_o[8]),
        .I2(load_i[1]),
        .O(\r_data[1]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__1 
       (.I0(writedata_i[17]),
        .I1(readdata_o[16]),
        .I2(load_i[2]),
        .O(\r_data[1]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__10 
       (.I0(writedata_i[89]),
        .I1(readdata_o[88]),
        .I2(load_i[11]),
        .O(\r_data[1]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__11 
       (.I0(writedata_i[97]),
        .I1(readdata_o[96]),
        .I2(load_i[12]),
        .O(\r_data[1]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair58" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__12 
       (.I0(writedata_i[105]),
        .I1(readdata_o[104]),
        .I2(load_i[13]),
        .O(\r_data[1]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair62" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__13 
       (.I0(writedata_i[113]),
        .I1(readdata_o[112]),
        .I2(load_i[14]),
        .O(\r_data[1]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair66" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__14 
       (.I0(writedata_i[121]),
        .I1(readdata_o[120]),
        .I2(load_i[15]),
        .O(\r_data[1]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair71" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__15 
       (.I0(writedata_i[129]),
        .I1(readdata_o[128]),
        .I2(load_i[16]),
        .O(\r_data[1]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair75" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__16 
       (.I0(writedata_i[137]),
        .I1(readdata_o[136]),
        .I2(load_i[17]),
        .O(\r_data[1]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair79" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__17 
       (.I0(writedata_i[145]),
        .I1(readdata_o[144]),
        .I2(load_i[18]),
        .O(\r_data[1]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair129" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__18 
       (.I0(writedata_i[153]),
        .I1(readdata_o[152]),
        .I2(load_i[19]),
        .O(\r_data[1]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__19 
       (.I0(writedata_i[161]),
        .I1(readdata_o[160]),
        .I2(load_i[20]),
        .O(\r_data[1]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__2 
       (.I0(writedata_i[25]),
        .I1(readdata_o[24]),
        .I2(load_i[3]),
        .O(\r_data[1]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair91" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__20 
       (.I0(writedata_i[169]),
        .I1(readdata_o[168]),
        .I2(load_i[21]),
        .O(\r_data[1]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair95" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__21 
       (.I0(writedata_i[177]),
        .I1(readdata_o[176]),
        .I2(load_i[22]),
        .O(\r_data[1]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair100" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__22 
       (.I0(writedata_i[185]),
        .I1(readdata_o[184]),
        .I2(load_i[23]),
        .O(\r_data[1]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair104" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__23 
       (.I0(writedata_i[193]),
        .I1(readdata_o[192]),
        .I2(load_i[24]),
        .O(\r_data[1]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair108" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__24 
       (.I0(writedata_i[201]),
        .I1(readdata_o[200]),
        .I2(load_i[25]),
        .O(\r_data[1]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair112" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__25 
       (.I0(writedata_i[209]),
        .I1(readdata_o[208]),
        .I2(load_i[26]),
        .O(\r_data[1]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair116" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__26 
       (.I0(writedata_i[217]),
        .I1(readdata_o[216]),
        .I2(load_i[27]),
        .O(\r_data[1]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair121" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__27 
       (.I0(writedata_i[225]),
        .I1(readdata_o[224]),
        .I2(load_i[28]),
        .O(\r_data[1]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__28 
       (.I0(writedata_i[233]),
        .I1(readdata_o[232]),
        .I2(load_i[29]),
        .O(\r_data[1]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair130" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__29 
       (.I0(writedata_i[241]),
        .I1(readdata_o[240]),
        .I2(load_i[30]),
        .O(\r_data[1]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__3 
       (.I0(writedata_i[33]),
        .I1(readdata_o[32]),
        .I2(load_i[4]),
        .O(\r_data[1]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair137" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__30 
       (.I0(writedata_i[249]),
        .I1(readdata_o[248]),
        .I2(load_i[31]),
        .O(\r_data[1]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__31 
       (.I0(writedata_i[257]),
        .I1(readdata_o[256]),
        .I2(load_i[32]),
        .O(\r_data[1]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair145" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__32 
       (.I0(writedata_i[265]),
        .I1(readdata_o[264]),
        .I2(load_i[33]),
        .O(\r_data[1]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair152" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__33 
       (.I0(writedata_i[273]),
        .I1(readdata_o[272]),
        .I2(load_i[34]),
        .O(\r_data[1]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair157" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__34 
       (.I0(writedata_i[281]),
        .I1(readdata_o[280]),
        .I2(load_i[35]),
        .O(\r_data[1]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair161" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__35 
       (.I0(writedata_i[289]),
        .I1(readdata_o[288]),
        .I2(load_i[36]),
        .O(\r_data[1]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair165" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__36 
       (.I0(writedata_i[297]),
        .I1(readdata_o[296]),
        .I2(load_i[37]),
        .O(\r_data[1]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair169" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__37 
       (.I0(writedata_i[305]),
        .I1(readdata_o[304]),
        .I2(load_i[38]),
        .O(\r_data[1]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair173" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__38 
       (.I0(writedata_i[313]),
        .I1(readdata_o[312]),
        .I2(load_i[39]),
        .O(\r_data[1]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair177" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__39 
       (.I0(writedata_i[321]),
        .I1(readdata_o[320]),
        .I2(load_i[40]),
        .O(\r_data[1]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__4 
       (.I0(writedata_i[41]),
        .I1(readdata_o[40]),
        .I2(load_i[5]),
        .O(\r_data[1]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair181" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__40 
       (.I0(writedata_i[329]),
        .I1(readdata_o[328]),
        .I2(load_i[41]),
        .O(\r_data[1]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair185" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__41 
       (.I0(writedata_i[337]),
        .I1(readdata_o[336]),
        .I2(load_i[42]),
        .O(\r_data[1]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair189" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__42 
       (.I0(writedata_i[345]),
        .I1(readdata_o[344]),
        .I2(load_i[43]),
        .O(\r_data[1]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair193" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__43 
       (.I0(writedata_i[353]),
        .I1(readdata_o[352]),
        .I2(load_i[44]),
        .O(\r_data[1]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair197" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__44 
       (.I0(writedata_i[361]),
        .I1(readdata_o[360]),
        .I2(load_i[45]),
        .O(\r_data[1]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair201" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__45 
       (.I0(writedata_i[369]),
        .I1(readdata_o[368]),
        .I2(load_i[46]),
        .O(\r_data[1]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair205" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__46 
       (.I0(writedata_i[377]),
        .I1(readdata_o[376]),
        .I2(load_i[47]),
        .O(\r_data[1]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair209" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__47 
       (.I0(writedata_i[385]),
        .I1(readdata_o[384]),
        .I2(load_i[48]),
        .O(\r_data[1]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__5 
       (.I0(writedata_i[49]),
        .I1(readdata_o[48]),
        .I2(load_i[6]),
        .O(\r_data[1]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__6 
       (.I0(writedata_i[57]),
        .I1(readdata_o[56]),
        .I2(load_i[7]),
        .O(\r_data[1]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__7 
       (.I0(writedata_i[65]),
        .I1(readdata_o[64]),
        .I2(load_i[8]),
        .O(\r_data[1]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__8 
       (.I0(writedata_i[73]),
        .I1(readdata_o[72]),
        .I2(load_i[9]),
        .O(\r_data[1]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[1]_i_1__9 
       (.I0(writedata_i[81]),
        .I1(readdata_o[80]),
        .I2(load_i[10]),
        .O(\r_data[1]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1 
       (.I0(writedata_i[2]),
        .I1(readdata_o[1]),
        .I2(load_i[0]),
        .O(\r_data[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__0 
       (.I0(writedata_i[10]),
        .I1(readdata_o[9]),
        .I2(load_i[1]),
        .O(\r_data[2]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__1 
       (.I0(writedata_i[18]),
        .I1(readdata_o[17]),
        .I2(load_i[2]),
        .O(\r_data[2]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair50" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__10 
       (.I0(writedata_i[90]),
        .I1(readdata_o[89]),
        .I2(load_i[11]),
        .O(\r_data[2]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair54" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__11 
       (.I0(writedata_i[98]),
        .I1(readdata_o[97]),
        .I2(load_i[12]),
        .O(\r_data[2]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__12 
       (.I0(writedata_i[106]),
        .I1(readdata_o[105]),
        .I2(load_i[13]),
        .O(\r_data[2]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__13 
       (.I0(writedata_i[114]),
        .I1(readdata_o[113]),
        .I2(load_i[14]),
        .O(\r_data[2]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__14 
       (.I0(writedata_i[122]),
        .I1(readdata_o[121]),
        .I2(load_i[15]),
        .O(\r_data[2]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__15 
       (.I0(writedata_i[130]),
        .I1(readdata_o[129]),
        .I2(load_i[16]),
        .O(\r_data[2]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__16 
       (.I0(writedata_i[138]),
        .I1(readdata_o[137]),
        .I2(load_i[17]),
        .O(\r_data[2]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__17 
       (.I0(writedata_i[146]),
        .I1(readdata_o[145]),
        .I2(load_i[18]),
        .O(\r_data[2]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__18 
       (.I0(writedata_i[154]),
        .I1(readdata_o[153]),
        .I2(load_i[19]),
        .O(\r_data[2]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__19 
       (.I0(writedata_i[162]),
        .I1(readdata_o[161]),
        .I2(load_i[20]),
        .O(\r_data[2]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__2 
       (.I0(writedata_i[26]),
        .I1(readdata_o[25]),
        .I2(load_i[3]),
        .O(\r_data[2]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__20 
       (.I0(writedata_i[170]),
        .I1(readdata_o[169]),
        .I2(load_i[21]),
        .O(\r_data[2]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__21 
       (.I0(writedata_i[178]),
        .I1(readdata_o[177]),
        .I2(load_i[22]),
        .O(\r_data[2]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__22 
       (.I0(writedata_i[186]),
        .I1(readdata_o[185]),
        .I2(load_i[23]),
        .O(\r_data[2]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__23 
       (.I0(writedata_i[194]),
        .I1(readdata_o[193]),
        .I2(load_i[24]),
        .O(\r_data[2]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__24 
       (.I0(writedata_i[202]),
        .I1(readdata_o[201]),
        .I2(load_i[25]),
        .O(\r_data[2]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__25 
       (.I0(writedata_i[210]),
        .I1(readdata_o[209]),
        .I2(load_i[26]),
        .O(\r_data[2]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__26 
       (.I0(writedata_i[218]),
        .I1(readdata_o[217]),
        .I2(load_i[27]),
        .O(\r_data[2]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__27 
       (.I0(writedata_i[226]),
        .I1(readdata_o[225]),
        .I2(load_i[28]),
        .O(\r_data[2]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair127" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__28 
       (.I0(writedata_i[234]),
        .I1(readdata_o[233]),
        .I2(load_i[29]),
        .O(\r_data[2]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__29 
       (.I0(writedata_i[242]),
        .I1(readdata_o[241]),
        .I2(load_i[30]),
        .O(\r_data[2]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__3 
       (.I0(writedata_i[34]),
        .I1(readdata_o[33]),
        .I2(load_i[4]),
        .O(\r_data[2]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__30 
       (.I0(writedata_i[250]),
        .I1(readdata_o[249]),
        .I2(load_i[31]),
        .O(\r_data[2]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair143" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__31 
       (.I0(writedata_i[258]),
        .I1(readdata_o[257]),
        .I2(load_i[32]),
        .O(\r_data[2]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__32 
       (.I0(writedata_i[266]),
        .I1(readdata_o[265]),
        .I2(load_i[33]),
        .O(\r_data[2]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__33 
       (.I0(writedata_i[274]),
        .I1(readdata_o[273]),
        .I2(load_i[34]),
        .O(\r_data[2]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__34 
       (.I0(writedata_i[282]),
        .I1(readdata_o[281]),
        .I2(load_i[35]),
        .O(\r_data[2]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__35 
       (.I0(writedata_i[290]),
        .I1(readdata_o[289]),
        .I2(load_i[36]),
        .O(\r_data[2]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__36 
       (.I0(writedata_i[298]),
        .I1(readdata_o[297]),
        .I2(load_i[37]),
        .O(\r_data[2]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__37 
       (.I0(writedata_i[306]),
        .I1(readdata_o[305]),
        .I2(load_i[38]),
        .O(\r_data[2]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__38 
       (.I0(writedata_i[314]),
        .I1(readdata_o[313]),
        .I2(load_i[39]),
        .O(\r_data[2]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__39 
       (.I0(writedata_i[322]),
        .I1(readdata_o[321]),
        .I2(load_i[40]),
        .O(\r_data[2]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__4 
       (.I0(writedata_i[42]),
        .I1(readdata_o[41]),
        .I2(load_i[5]),
        .O(\r_data[2]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__40 
       (.I0(writedata_i[330]),
        .I1(readdata_o[329]),
        .I2(load_i[41]),
        .O(\r_data[2]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__41 
       (.I0(writedata_i[338]),
        .I1(readdata_o[337]),
        .I2(load_i[42]),
        .O(\r_data[2]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__42 
       (.I0(writedata_i[346]),
        .I1(readdata_o[345]),
        .I2(load_i[43]),
        .O(\r_data[2]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__43 
       (.I0(writedata_i[354]),
        .I1(readdata_o[353]),
        .I2(load_i[44]),
        .O(\r_data[2]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__44 
       (.I0(writedata_i[362]),
        .I1(readdata_o[361]),
        .I2(load_i[45]),
        .O(\r_data[2]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__45 
       (.I0(writedata_i[370]),
        .I1(readdata_o[369]),
        .I2(load_i[46]),
        .O(\r_data[2]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__46 
       (.I0(writedata_i[378]),
        .I1(readdata_o[377]),
        .I2(load_i[47]),
        .O(\r_data[2]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__47 
       (.I0(writedata_i[386]),
        .I1(readdata_o[385]),
        .I2(load_i[48]),
        .O(\r_data[2]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__5 
       (.I0(writedata_i[50]),
        .I1(readdata_o[49]),
        .I2(load_i[6]),
        .O(\r_data[2]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__6 
       (.I0(writedata_i[58]),
        .I1(readdata_o[57]),
        .I2(load_i[7]),
        .O(\r_data[2]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__7 
       (.I0(writedata_i[66]),
        .I1(readdata_o[65]),
        .I2(load_i[8]),
        .O(\r_data[2]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__8 
       (.I0(writedata_i[74]),
        .I1(readdata_o[73]),
        .I2(load_i[9]),
        .O(\r_data[2]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[2]_i_1__9 
       (.I0(writedata_i[82]),
        .I1(readdata_o[81]),
        .I2(load_i[10]),
        .O(\r_data[2]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1 
       (.I0(writedata_i[3]),
        .I1(readdata_o[2]),
        .I2(load_i[0]),
        .O(\r_data[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__0 
       (.I0(writedata_i[11]),
        .I1(readdata_o[10]),
        .I2(load_i[1]),
        .O(\r_data[3]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__1 
       (.I0(writedata_i[19]),
        .I1(readdata_o[18]),
        .I2(load_i[2]),
        .O(\r_data[3]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair51" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__10 
       (.I0(writedata_i[91]),
        .I1(readdata_o[90]),
        .I2(load_i[11]),
        .O(\r_data[3]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair55" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__11 
       (.I0(writedata_i[99]),
        .I1(readdata_o[98]),
        .I2(load_i[12]),
        .O(\r_data[3]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair59" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__12 
       (.I0(writedata_i[107]),
        .I1(readdata_o[106]),
        .I2(load_i[13]),
        .O(\r_data[3]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair63" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__13 
       (.I0(writedata_i[115]),
        .I1(readdata_o[114]),
        .I2(load_i[14]),
        .O(\r_data[3]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair67" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__14 
       (.I0(writedata_i[123]),
        .I1(readdata_o[122]),
        .I2(load_i[15]),
        .O(\r_data[3]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair72" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__15 
       (.I0(writedata_i[131]),
        .I1(readdata_o[130]),
        .I2(load_i[16]),
        .O(\r_data[3]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair76" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__16 
       (.I0(writedata_i[139]),
        .I1(readdata_o[138]),
        .I2(load_i[17]),
        .O(\r_data[3]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair98" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__17 
       (.I0(writedata_i[147]),
        .I1(readdata_o[146]),
        .I2(load_i[18]),
        .O(\r_data[3]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair134" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__18 
       (.I0(writedata_i[155]),
        .I1(readdata_o[154]),
        .I2(load_i[19]),
        .O(\r_data[3]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair149" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__19 
       (.I0(writedata_i[163]),
        .I1(readdata_o[162]),
        .I2(load_i[20]),
        .O(\r_data[3]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__2 
       (.I0(writedata_i[27]),
        .I1(readdata_o[26]),
        .I2(load_i[3]),
        .O(\r_data[3]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair92" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__20 
       (.I0(writedata_i[171]),
        .I1(readdata_o[170]),
        .I2(load_i[21]),
        .O(\r_data[3]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair96" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__21 
       (.I0(writedata_i[179]),
        .I1(readdata_o[178]),
        .I2(load_i[22]),
        .O(\r_data[3]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair101" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__22 
       (.I0(writedata_i[187]),
        .I1(readdata_o[186]),
        .I2(load_i[23]),
        .O(\r_data[3]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair105" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__23 
       (.I0(writedata_i[195]),
        .I1(readdata_o[194]),
        .I2(load_i[24]),
        .O(\r_data[3]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair109" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__24 
       (.I0(writedata_i[203]),
        .I1(readdata_o[202]),
        .I2(load_i[25]),
        .O(\r_data[3]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair113" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__25 
       (.I0(writedata_i[211]),
        .I1(readdata_o[210]),
        .I2(load_i[26]),
        .O(\r_data[3]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair117" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__26 
       (.I0(writedata_i[219]),
        .I1(readdata_o[218]),
        .I2(load_i[27]),
        .O(\r_data[3]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__27 
       (.I0(writedata_i[227]),
        .I1(readdata_o[226]),
        .I2(load_i[28]),
        .O(\r_data[3]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__28 
       (.I0(writedata_i[235]),
        .I1(readdata_o[234]),
        .I2(load_i[29]),
        .O(\r_data[3]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair132" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__29 
       (.I0(writedata_i[243]),
        .I1(readdata_o[242]),
        .I2(load_i[30]),
        .O(\r_data[3]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__3 
       (.I0(writedata_i[35]),
        .I1(readdata_o[34]),
        .I2(load_i[4]),
        .O(\r_data[3]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__30 
       (.I0(writedata_i[251]),
        .I1(readdata_o[250]),
        .I2(load_i[31]),
        .O(\r_data[3]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__31 
       (.I0(writedata_i[259]),
        .I1(readdata_o[258]),
        .I2(load_i[32]),
        .O(\r_data[3]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair147" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__32 
       (.I0(writedata_i[267]),
        .I1(readdata_o[266]),
        .I2(load_i[33]),
        .O(\r_data[3]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__33 
       (.I0(writedata_i[275]),
        .I1(readdata_o[274]),
        .I2(load_i[34]),
        .O(\r_data[3]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair158" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__34 
       (.I0(writedata_i[283]),
        .I1(readdata_o[282]),
        .I2(load_i[35]),
        .O(\r_data[3]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair162" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__35 
       (.I0(writedata_i[291]),
        .I1(readdata_o[290]),
        .I2(load_i[36]),
        .O(\r_data[3]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair166" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__36 
       (.I0(writedata_i[299]),
        .I1(readdata_o[298]),
        .I2(load_i[37]),
        .O(\r_data[3]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair170" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__37 
       (.I0(writedata_i[307]),
        .I1(readdata_o[306]),
        .I2(load_i[38]),
        .O(\r_data[3]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair174" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__38 
       (.I0(writedata_i[315]),
        .I1(readdata_o[314]),
        .I2(load_i[39]),
        .O(\r_data[3]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair178" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__39 
       (.I0(writedata_i[323]),
        .I1(readdata_o[322]),
        .I2(load_i[40]),
        .O(\r_data[3]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__4 
       (.I0(writedata_i[43]),
        .I1(readdata_o[42]),
        .I2(load_i[5]),
        .O(\r_data[3]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair182" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__40 
       (.I0(writedata_i[331]),
        .I1(readdata_o[330]),
        .I2(load_i[41]),
        .O(\r_data[3]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair186" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__41 
       (.I0(writedata_i[339]),
        .I1(readdata_o[338]),
        .I2(load_i[42]),
        .O(\r_data[3]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair190" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__42 
       (.I0(writedata_i[347]),
        .I1(readdata_o[346]),
        .I2(load_i[43]),
        .O(\r_data[3]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair194" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__43 
       (.I0(writedata_i[355]),
        .I1(readdata_o[354]),
        .I2(load_i[44]),
        .O(\r_data[3]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair198" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__44 
       (.I0(writedata_i[363]),
        .I1(readdata_o[362]),
        .I2(load_i[45]),
        .O(\r_data[3]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair202" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__45 
       (.I0(writedata_i[371]),
        .I1(readdata_o[370]),
        .I2(load_i[46]),
        .O(\r_data[3]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair206" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__46 
       (.I0(writedata_i[379]),
        .I1(readdata_o[378]),
        .I2(load_i[47]),
        .O(\r_data[3]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair210" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__47 
       (.I0(writedata_i[387]),
        .I1(readdata_o[386]),
        .I2(load_i[48]),
        .O(\r_data[3]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__5 
       (.I0(writedata_i[51]),
        .I1(readdata_o[50]),
        .I2(load_i[6]),
        .O(\r_data[3]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__6 
       (.I0(writedata_i[59]),
        .I1(readdata_o[58]),
        .I2(load_i[7]),
        .O(\r_data[3]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__7 
       (.I0(writedata_i[67]),
        .I1(readdata_o[66]),
        .I2(load_i[8]),
        .O(\r_data[3]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__8 
       (.I0(writedata_i[75]),
        .I1(readdata_o[74]),
        .I2(load_i[9]),
        .O(\r_data[3]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[3]_i_1__9 
       (.I0(writedata_i[83]),
        .I1(readdata_o[82]),
        .I2(load_i[10]),
        .O(\r_data[3]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair293" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1 
       (.I0(writedata_i[4]),
        .I1(readdata_o[3]),
        .I2(load_i[0]),
        .O(\r_data[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair289" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__0 
       (.I0(writedata_i[12]),
        .I1(readdata_o[11]),
        .I2(load_i[1]),
        .O(\r_data[4]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair285" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__1 
       (.I0(writedata_i[20]),
        .I1(readdata_o[19]),
        .I2(load_i[2]),
        .O(\r_data[4]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__10 
       (.I0(writedata_i[92]),
        .I1(readdata_o[91]),
        .I2(load_i[11]),
        .O(\r_data[4]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__11 
       (.I0(writedata_i[100]),
        .I1(readdata_o[99]),
        .I2(load_i[12]),
        .O(\r_data[4]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__12 
       (.I0(writedata_i[108]),
        .I1(readdata_o[107]),
        .I2(load_i[13]),
        .O(\r_data[4]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__13 
       (.I0(writedata_i[116]),
        .I1(readdata_o[115]),
        .I2(load_i[14]),
        .O(\r_data[4]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__14 
       (.I0(writedata_i[124]),
        .I1(readdata_o[123]),
        .I2(load_i[15]),
        .O(\r_data[4]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__15 
       (.I0(writedata_i[132]),
        .I1(readdata_o[131]),
        .I2(load_i[16]),
        .O(\r_data[4]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__16 
       (.I0(writedata_i[140]),
        .I1(readdata_o[139]),
        .I2(load_i[17]),
        .O(\r_data[4]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__17 
       (.I0(writedata_i[148]),
        .I1(readdata_o[147]),
        .I2(load_i[18]),
        .O(\r_data[4]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__18 
       (.I0(writedata_i[156]),
        .I1(readdata_o[155]),
        .I2(load_i[19]),
        .O(\r_data[4]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__19 
       (.I0(writedata_i[164]),
        .I1(readdata_o[163]),
        .I2(load_i[20]),
        .O(\r_data[4]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair281" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__2 
       (.I0(writedata_i[28]),
        .I1(readdata_o[27]),
        .I2(load_i[3]),
        .O(\r_data[4]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__20 
       (.I0(writedata_i[172]),
        .I1(readdata_o[171]),
        .I2(load_i[21]),
        .O(\r_data[4]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__21 
       (.I0(writedata_i[180]),
        .I1(readdata_o[179]),
        .I2(load_i[22]),
        .O(\r_data[4]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__22 
       (.I0(writedata_i[188]),
        .I1(readdata_o[187]),
        .I2(load_i[23]),
        .O(\r_data[4]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__23 
       (.I0(writedata_i[196]),
        .I1(readdata_o[195]),
        .I2(load_i[24]),
        .O(\r_data[4]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__24 
       (.I0(writedata_i[204]),
        .I1(readdata_o[203]),
        .I2(load_i[25]),
        .O(\r_data[4]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__25 
       (.I0(writedata_i[212]),
        .I1(readdata_o[211]),
        .I2(load_i[26]),
        .O(\r_data[4]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__26 
       (.I0(writedata_i[220]),
        .I1(readdata_o[219]),
        .I2(load_i[27]),
        .O(\r_data[4]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair124" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__27 
       (.I0(writedata_i[228]),
        .I1(readdata_o[227]),
        .I2(load_i[28]),
        .O(\r_data[4]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair223" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__28 
       (.I0(writedata_i[236]),
        .I1(readdata_o[235]),
        .I2(load_i[29]),
        .O(\r_data[4]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__29 
       (.I0(writedata_i[244]),
        .I1(readdata_o[243]),
        .I2(load_i[30]),
        .O(\r_data[4]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair277" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__3 
       (.I0(writedata_i[36]),
        .I1(readdata_o[35]),
        .I2(load_i[4]),
        .O(\r_data[4]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair140" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__30 
       (.I0(writedata_i[252]),
        .I1(readdata_o[251]),
        .I2(load_i[31]),
        .O(\r_data[4]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair243" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__31 
       (.I0(writedata_i[260]),
        .I1(readdata_o[259]),
        .I2(load_i[32]),
        .O(\r_data[4]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__32 
       (.I0(writedata_i[268]),
        .I1(readdata_o[267]),
        .I2(load_i[33]),
        .O(\r_data[4]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair155" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__33 
       (.I0(writedata_i[276]),
        .I1(readdata_o[275]),
        .I2(load_i[34]),
        .O(\r_data[4]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__34 
       (.I0(writedata_i[284]),
        .I1(readdata_o[283]),
        .I2(load_i[35]),
        .O(\r_data[4]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__35 
       (.I0(writedata_i[292]),
        .I1(readdata_o[291]),
        .I2(load_i[36]),
        .O(\r_data[4]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__36 
       (.I0(writedata_i[300]),
        .I1(readdata_o[299]),
        .I2(load_i[37]),
        .O(\r_data[4]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__37 
       (.I0(writedata_i[308]),
        .I1(readdata_o[307]),
        .I2(load_i[38]),
        .O(\r_data[4]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__38 
       (.I0(writedata_i[316]),
        .I1(readdata_o[315]),
        .I2(load_i[39]),
        .O(\r_data[4]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__39 
       (.I0(writedata_i[324]),
        .I1(readdata_o[323]),
        .I2(load_i[40]),
        .O(\r_data[4]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair270" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__4 
       (.I0(writedata_i[44]),
        .I1(readdata_o[43]),
        .I2(load_i[5]),
        .O(\r_data[4]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__40 
       (.I0(writedata_i[332]),
        .I1(readdata_o[331]),
        .I2(load_i[41]),
        .O(\r_data[4]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__41 
       (.I0(writedata_i[340]),
        .I1(readdata_o[339]),
        .I2(load_i[42]),
        .O(\r_data[4]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__42 
       (.I0(writedata_i[348]),
        .I1(readdata_o[347]),
        .I2(load_i[43]),
        .O(\r_data[4]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__43 
       (.I0(writedata_i[356]),
        .I1(readdata_o[355]),
        .I2(load_i[44]),
        .O(\r_data[4]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__44 
       (.I0(writedata_i[364]),
        .I1(readdata_o[363]),
        .I2(load_i[45]),
        .O(\r_data[4]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__45 
       (.I0(writedata_i[372]),
        .I1(readdata_o[371]),
        .I2(load_i[46]),
        .O(\r_data[4]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__46 
       (.I0(writedata_i[380]),
        .I1(readdata_o[379]),
        .I2(load_i[47]),
        .O(\r_data[4]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__47 
       (.I0(writedata_i[388]),
        .I1(readdata_o[387]),
        .I2(load_i[48]),
        .O(\r_data[4]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair153" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__5 
       (.I0(writedata_i[52]),
        .I1(readdata_o[51]),
        .I2(load_i[6]),
        .O(\r_data[4]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair138" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__6 
       (.I0(writedata_i[60]),
        .I1(readdata_o[59]),
        .I2(load_i[7]),
        .O(\r_data[4]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair122" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__7 
       (.I0(writedata_i[68]),
        .I1(readdata_o[67]),
        .I2(load_i[8]),
        .O(\r_data[4]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair87" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__8 
       (.I0(writedata_i[76]),
        .I1(readdata_o[75]),
        .I2(load_i[9]),
        .O(\r_data[4]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair83" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[4]_i_1__9 
       (.I0(writedata_i[84]),
        .I1(readdata_o[83]),
        .I2(load_i[10]),
        .O(\r_data[4]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair292" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1 
       (.I0(writedata_i[5]),
        .I1(readdata_o[4]),
        .I2(load_i[0]),
        .O(\r_data[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair288" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__0 
       (.I0(writedata_i[13]),
        .I1(readdata_o[12]),
        .I2(load_i[1]),
        .O(\r_data[5]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair284" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__1 
       (.I0(writedata_i[21]),
        .I1(readdata_o[20]),
        .I2(load_i[2]),
        .O(\r_data[5]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair52" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__10 
       (.I0(writedata_i[93]),
        .I1(readdata_o[92]),
        .I2(load_i[11]),
        .O(\r_data[5]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair56" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__11 
       (.I0(writedata_i[101]),
        .I1(readdata_o[100]),
        .I2(load_i[12]),
        .O(\r_data[5]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair60" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__12 
       (.I0(writedata_i[109]),
        .I1(readdata_o[108]),
        .I2(load_i[13]),
        .O(\r_data[5]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair64" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__13 
       (.I0(writedata_i[117]),
        .I1(readdata_o[116]),
        .I2(load_i[14]),
        .O(\r_data[5]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair68" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__14 
       (.I0(writedata_i[125]),
        .I1(readdata_o[124]),
        .I2(load_i[15]),
        .O(\r_data[5]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair73" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__15 
       (.I0(writedata_i[133]),
        .I1(readdata_o[132]),
        .I2(load_i[16]),
        .O(\r_data[5]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair77" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__16 
       (.I0(writedata_i[141]),
        .I1(readdata_o[140]),
        .I2(load_i[17]),
        .O(\r_data[5]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair123" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__17 
       (.I0(writedata_i[149]),
        .I1(readdata_o[148]),
        .I2(load_i[18]),
        .O(\r_data[5]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair139" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__18 
       (.I0(writedata_i[157]),
        .I1(readdata_o[156]),
        .I2(load_i[19]),
        .O(\r_data[5]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair89" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__19 
       (.I0(writedata_i[165]),
        .I1(readdata_o[164]),
        .I2(load_i[20]),
        .O(\r_data[5]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair280" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__2 
       (.I0(writedata_i[29]),
        .I1(readdata_o[28]),
        .I2(load_i[3]),
        .O(\r_data[5]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair93" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__20 
       (.I0(writedata_i[173]),
        .I1(readdata_o[172]),
        .I2(load_i[21]),
        .O(\r_data[5]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair97" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__21 
       (.I0(writedata_i[181]),
        .I1(readdata_o[180]),
        .I2(load_i[22]),
        .O(\r_data[5]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair102" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__22 
       (.I0(writedata_i[189]),
        .I1(readdata_o[188]),
        .I2(load_i[23]),
        .O(\r_data[5]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair106" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__23 
       (.I0(writedata_i[197]),
        .I1(readdata_o[196]),
        .I2(load_i[24]),
        .O(\r_data[5]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair110" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__24 
       (.I0(writedata_i[205]),
        .I1(readdata_o[204]),
        .I2(load_i[25]),
        .O(\r_data[5]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair114" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__25 
       (.I0(writedata_i[213]),
        .I1(readdata_o[212]),
        .I2(load_i[26]),
        .O(\r_data[5]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair118" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__26 
       (.I0(writedata_i[221]),
        .I1(readdata_o[220]),
        .I2(load_i[27]),
        .O(\r_data[5]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__27 
       (.I0(writedata_i[229]),
        .I1(readdata_o[228]),
        .I2(load_i[28]),
        .O(\r_data[5]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair128" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__28 
       (.I0(writedata_i[237]),
        .I1(readdata_o[236]),
        .I2(load_i[29]),
        .O(\r_data[5]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__29 
       (.I0(writedata_i[245]),
        .I1(readdata_o[244]),
        .I2(load_i[30]),
        .O(\r_data[5]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair276" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__3 
       (.I0(writedata_i[37]),
        .I1(readdata_o[36]),
        .I2(load_i[4]),
        .O(\r_data[5]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__30 
       (.I0(writedata_i[253]),
        .I1(readdata_o[252]),
        .I2(load_i[31]),
        .O(\r_data[5]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair144" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__31 
       (.I0(writedata_i[261]),
        .I1(readdata_o[260]),
        .I2(load_i[32]),
        .O(\r_data[5]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__32 
       (.I0(writedata_i[269]),
        .I1(readdata_o[268]),
        .I2(load_i[33]),
        .O(\r_data[5]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__33 
       (.I0(writedata_i[277]),
        .I1(readdata_o[276]),
        .I2(load_i[34]),
        .O(\r_data[5]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair159" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__34 
       (.I0(writedata_i[285]),
        .I1(readdata_o[284]),
        .I2(load_i[35]),
        .O(\r_data[5]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair163" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__35 
       (.I0(writedata_i[293]),
        .I1(readdata_o[292]),
        .I2(load_i[36]),
        .O(\r_data[5]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair167" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__36 
       (.I0(writedata_i[301]),
        .I1(readdata_o[300]),
        .I2(load_i[37]),
        .O(\r_data[5]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair171" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__37 
       (.I0(writedata_i[309]),
        .I1(readdata_o[308]),
        .I2(load_i[38]),
        .O(\r_data[5]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair175" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__38 
       (.I0(writedata_i[317]),
        .I1(readdata_o[316]),
        .I2(load_i[39]),
        .O(\r_data[5]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair179" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__39 
       (.I0(writedata_i[325]),
        .I1(readdata_o[324]),
        .I2(load_i[40]),
        .O(\r_data[5]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair268" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__4 
       (.I0(writedata_i[45]),
        .I1(readdata_o[44]),
        .I2(load_i[5]),
        .O(\r_data[5]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair183" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__40 
       (.I0(writedata_i[333]),
        .I1(readdata_o[332]),
        .I2(load_i[41]),
        .O(\r_data[5]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair187" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__41 
       (.I0(writedata_i[341]),
        .I1(readdata_o[340]),
        .I2(load_i[42]),
        .O(\r_data[5]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair191" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__42 
       (.I0(writedata_i[349]),
        .I1(readdata_o[348]),
        .I2(load_i[43]),
        .O(\r_data[5]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair195" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__43 
       (.I0(writedata_i[357]),
        .I1(readdata_o[356]),
        .I2(load_i[44]),
        .O(\r_data[5]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair199" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__44 
       (.I0(writedata_i[365]),
        .I1(readdata_o[364]),
        .I2(load_i[45]),
        .O(\r_data[5]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair203" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__45 
       (.I0(writedata_i[373]),
        .I1(readdata_o[372]),
        .I2(load_i[46]),
        .O(\r_data[5]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair207" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__46 
       (.I0(writedata_i[381]),
        .I1(readdata_o[380]),
        .I2(load_i[47]),
        .O(\r_data[5]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair211" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__47 
       (.I0(writedata_i[389]),
        .I1(readdata_o[388]),
        .I2(load_i[48]),
        .O(\r_data[5]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair151" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__5 
       (.I0(writedata_i[53]),
        .I1(readdata_o[52]),
        .I2(load_i[6]),
        .O(\r_data[5]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair136" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__6 
       (.I0(writedata_i[61]),
        .I1(readdata_o[60]),
        .I2(load_i[7]),
        .O(\r_data[5]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair120" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__7 
       (.I0(writedata_i[69]),
        .I1(readdata_o[68]),
        .I2(load_i[8]),
        .O(\r_data[5]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair86" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__8 
       (.I0(writedata_i[77]),
        .I1(readdata_o[76]),
        .I2(load_i[9]),
        .O(\r_data[5]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair82" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[5]_i_1__9 
       (.I0(writedata_i[85]),
        .I1(readdata_o[84]),
        .I2(load_i[10]),
        .O(\r_data[5]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair291" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1 
       (.I0(writedata_i[6]),
        .I1(readdata_o[5]),
        .I2(load_i[0]),
        .O(\r_data[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair287" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__0 
       (.I0(writedata_i[14]),
        .I1(readdata_o[13]),
        .I2(load_i[1]),
        .O(\r_data[6]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair283" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__1 
       (.I0(writedata_i[22]),
        .I1(readdata_o[21]),
        .I2(load_i[2]),
        .O(\r_data[6]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__10 
       (.I0(writedata_i[94]),
        .I1(readdata_o[93]),
        .I2(load_i[11]),
        .O(\r_data[6]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__11 
       (.I0(writedata_i[102]),
        .I1(readdata_o[101]),
        .I2(load_i[12]),
        .O(\r_data[6]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__12 
       (.I0(writedata_i[110]),
        .I1(readdata_o[109]),
        .I2(load_i[13]),
        .O(\r_data[6]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__13 
       (.I0(writedata_i[118]),
        .I1(readdata_o[117]),
        .I2(load_i[14]),
        .O(\r_data[6]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__14 
       (.I0(writedata_i[126]),
        .I1(readdata_o[125]),
        .I2(load_i[15]),
        .O(\r_data[6]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__15 
       (.I0(writedata_i[134]),
        .I1(readdata_o[133]),
        .I2(load_i[16]),
        .O(\r_data[6]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__16 
       (.I0(writedata_i[142]),
        .I1(readdata_o[141]),
        .I2(load_i[17]),
        .O(\r_data[6]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__17 
       (.I0(writedata_i[150]),
        .I1(readdata_o[149]),
        .I2(load_i[18]),
        .O(\r_data[6]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__18 
       (.I0(writedata_i[158]),
        .I1(readdata_o[157]),
        .I2(load_i[19]),
        .O(\r_data[6]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair154" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__19 
       (.I0(writedata_i[166]),
        .I1(readdata_o[165]),
        .I2(load_i[20]),
        .O(\r_data[6]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair279" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__2 
       (.I0(writedata_i[30]),
        .I1(readdata_o[29]),
        .I2(load_i[3]),
        .O(\r_data[6]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__20 
       (.I0(writedata_i[174]),
        .I1(readdata_o[173]),
        .I2(load_i[21]),
        .O(\r_data[6]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__21 
       (.I0(writedata_i[182]),
        .I1(readdata_o[181]),
        .I2(load_i[22]),
        .O(\r_data[6]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__22 
       (.I0(writedata_i[190]),
        .I1(readdata_o[189]),
        .I2(load_i[23]),
        .O(\r_data[6]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__23 
       (.I0(writedata_i[198]),
        .I1(readdata_o[197]),
        .I2(load_i[24]),
        .O(\r_data[6]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__24 
       (.I0(writedata_i[206]),
        .I1(readdata_o[205]),
        .I2(load_i[25]),
        .O(\r_data[6]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__25 
       (.I0(writedata_i[214]),
        .I1(readdata_o[213]),
        .I2(load_i[26]),
        .O(\r_data[6]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__26 
       (.I0(writedata_i[222]),
        .I1(readdata_o[221]),
        .I2(load_i[27]),
        .O(\r_data[6]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair218" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__27 
       (.I0(writedata_i[230]),
        .I1(readdata_o[229]),
        .I2(load_i[28]),
        .O(\r_data[6]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__28 
       (.I0(writedata_i[238]),
        .I1(readdata_o[237]),
        .I2(load_i[29]),
        .O(\r_data[6]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair135" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__29 
       (.I0(writedata_i[246]),
        .I1(readdata_o[245]),
        .I2(load_i[30]),
        .O(\r_data[6]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair275" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__3 
       (.I0(writedata_i[38]),
        .I1(readdata_o[37]),
        .I2(load_i[4]),
        .O(\r_data[6]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair238" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__30 
       (.I0(writedata_i[254]),
        .I1(readdata_o[253]),
        .I2(load_i[31]),
        .O(\r_data[6]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__31 
       (.I0(writedata_i[262]),
        .I1(readdata_o[261]),
        .I2(load_i[32]),
        .O(\r_data[6]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair150" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__32 
       (.I0(writedata_i[270]),
        .I1(readdata_o[269]),
        .I2(load_i[33]),
        .O(\r_data[6]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair258" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__33 
       (.I0(writedata_i[278]),
        .I1(readdata_o[277]),
        .I2(load_i[34]),
        .O(\r_data[6]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__34 
       (.I0(writedata_i[286]),
        .I1(readdata_o[285]),
        .I2(load_i[35]),
        .O(\r_data[6]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__35 
       (.I0(writedata_i[294]),
        .I1(readdata_o[293]),
        .I2(load_i[36]),
        .O(\r_data[6]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__36 
       (.I0(writedata_i[302]),
        .I1(readdata_o[301]),
        .I2(load_i[37]),
        .O(\r_data[6]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__37 
       (.I0(writedata_i[310]),
        .I1(readdata_o[309]),
        .I2(load_i[38]),
        .O(\r_data[6]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__38 
       (.I0(writedata_i[318]),
        .I1(readdata_o[317]),
        .I2(load_i[39]),
        .O(\r_data[6]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__39 
       (.I0(writedata_i[326]),
        .I1(readdata_o[325]),
        .I2(load_i[40]),
        .O(\r_data[6]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair266" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__4 
       (.I0(writedata_i[46]),
        .I1(readdata_o[45]),
        .I2(load_i[5]),
        .O(\r_data[6]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__40 
       (.I0(writedata_i[334]),
        .I1(readdata_o[333]),
        .I2(load_i[41]),
        .O(\r_data[6]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__41 
       (.I0(writedata_i[342]),
        .I1(readdata_o[341]),
        .I2(load_i[42]),
        .O(\r_data[6]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__42 
       (.I0(writedata_i[350]),
        .I1(readdata_o[349]),
        .I2(load_i[43]),
        .O(\r_data[6]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__43 
       (.I0(writedata_i[358]),
        .I1(readdata_o[357]),
        .I2(load_i[44]),
        .O(\r_data[6]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__44 
       (.I0(writedata_i[366]),
        .I1(readdata_o[365]),
        .I2(load_i[45]),
        .O(\r_data[6]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__45 
       (.I0(writedata_i[374]),
        .I1(readdata_o[373]),
        .I2(load_i[46]),
        .O(\r_data[6]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__46 
       (.I0(writedata_i[382]),
        .I1(readdata_o[381]),
        .I2(load_i[47]),
        .O(\r_data[6]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__47 
       (.I0(writedata_i[390]),
        .I1(readdata_o[389]),
        .I2(load_i[48]),
        .O(\r_data[6]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair148" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__5 
       (.I0(writedata_i[54]),
        .I1(readdata_o[53]),
        .I2(load_i[6]),
        .O(\r_data[6]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair133" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__6 
       (.I0(writedata_i[62]),
        .I1(readdata_o[61]),
        .I2(load_i[7]),
        .O(\r_data[6]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair69" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__7 
       (.I0(writedata_i[70]),
        .I1(readdata_o[69]),
        .I2(load_i[8]),
        .O(\r_data[6]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair85" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__8 
       (.I0(writedata_i[78]),
        .I1(readdata_o[77]),
        .I2(load_i[9]),
        .O(\r_data[6]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair81" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[6]_i_1__9 
       (.I0(writedata_i[86]),
        .I1(readdata_o[85]),
        .I2(load_i[10]),
        .O(\r_data[6]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1 
       (.I0(load_i[0]),
        .I1(w_run_up_2),
        .I2(w_run),
        .O(\r_data[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__0 
       (.I0(load_i[1]),
        .I1(w_run_up_3),
        .I2(w_run_up_1),
        .O(\r_data[7]_i_1__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__1 
       (.I0(load_i[2]),
        .I1(w_run_up_4),
        .I2(w_run_up_2),
        .O(\r_data[7]_i_1__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__10 
       (.I0(load_i[11]),
        .I1(w_run_up_13),
        .I2(w_run_up_11),
        .O(\r_data[7]_i_1__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__11 
       (.I0(load_i[12]),
        .I1(w_run_up_14),
        .I2(w_run_up_12),
        .O(\r_data[7]_i_1__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__12 
       (.I0(load_i[13]),
        .I1(w_run_up_15),
        .I2(w_run_up_13),
        .O(\r_data[7]_i_1__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__13 
       (.I0(load_i[14]),
        .I1(w_run_up_16),
        .I2(w_run_up_14),
        .O(\r_data[7]_i_1__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__14 
       (.I0(load_i[15]),
        .I1(w_run_up_17),
        .I2(w_run_up_15),
        .O(\r_data[7]_i_1__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__15 
       (.I0(load_i[16]),
        .I1(w_run_up_18),
        .I2(w_run_up_16),
        .O(\r_data[7]_i_1__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__16 
       (.I0(load_i[17]),
        .I1(w_run_up_19),
        .I2(w_run_up_17),
        .O(\r_data[7]_i_1__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__17 
       (.I0(load_i[18]),
        .I1(w_run_up_20),
        .I2(w_run_up_18),
        .O(\r_data[7]_i_1__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__18 
       (.I0(load_i[19]),
        .I1(w_run_up_21),
        .I2(w_run_up_19),
        .O(\r_data[7]_i_1__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__19 
       (.I0(load_i[20]),
        .I1(w_run_up_22),
        .I2(w_run_up_20),
        .O(\r_data[7]_i_1__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__2 
       (.I0(load_i[3]),
        .I1(w_run_up_5),
        .I2(w_run_up_3),
        .O(\r_data[7]_i_1__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__20 
       (.I0(load_i[21]),
        .I1(w_run_up_23),
        .I2(w_run_up_21),
        .O(\r_data[7]_i_1__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__21 
       (.I0(load_i[22]),
        .I1(w_run_up_24),
        .I2(w_run_up_22),
        .O(\r_data[7]_i_1__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__22 
       (.I0(load_i[23]),
        .I1(w_run_up_25),
        .I2(w_run_up_23),
        .O(\r_data[7]_i_1__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__23 
       (.I0(load_i[24]),
        .I1(w_run_up_26),
        .I2(w_run_up_24),
        .O(\r_data[7]_i_1__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__24 
       (.I0(load_i[25]),
        .I1(w_run_up_27),
        .I2(w_run_up_25),
        .O(\r_data[7]_i_1__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__25 
       (.I0(load_i[26]),
        .I1(w_run_up_28),
        .I2(w_run_up_26),
        .O(\r_data[7]_i_1__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__26 
       (.I0(load_i[27]),
        .I1(w_run_up_29),
        .I2(w_run_up_27),
        .O(\r_data[7]_i_1__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__27 
       (.I0(load_i[28]),
        .I1(w_run_up_30),
        .I2(w_run_up_28),
        .O(\r_data[7]_i_1__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__28 
       (.I0(load_i[29]),
        .I1(w_run_up_31),
        .I2(w_run_up_29),
        .O(\r_data[7]_i_1__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__29 
       (.I0(load_i[30]),
        .I1(w_run_up_32),
        .I2(w_run_up_30),
        .O(\r_data[7]_i_1__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__3 
       (.I0(load_i[4]),
        .I1(w_run_up_6),
        .I2(w_run_up_4),
        .O(\r_data[7]_i_1__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__30 
       (.I0(load_i[31]),
        .I1(w_run_up_33),
        .I2(w_run_up_31),
        .O(\r_data[7]_i_1__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__31 
       (.I0(load_i[32]),
        .I1(w_run_up_34),
        .I2(w_run_up_32),
        .O(\r_data[7]_i_1__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__32 
       (.I0(load_i[33]),
        .I1(w_run_up_35),
        .I2(w_run_up_33),
        .O(\r_data[7]_i_1__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__33 
       (.I0(load_i[34]),
        .I1(w_run_up_36),
        .I2(w_run_up_34),
        .O(\r_data[7]_i_1__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__34 
       (.I0(load_i[35]),
        .I1(w_run_up_37),
        .I2(w_run_up_35),
        .O(\r_data[7]_i_1__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__35 
       (.I0(load_i[36]),
        .I1(w_run_up_38),
        .I2(w_run_up_36),
        .O(\r_data[7]_i_1__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__36 
       (.I0(load_i[37]),
        .I1(w_run_up_39),
        .I2(w_run_up_37),
        .O(\r_data[7]_i_1__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__37 
       (.I0(load_i[38]),
        .I1(w_run_up_40),
        .I2(w_run_up_38),
        .O(\r_data[7]_i_1__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__38 
       (.I0(load_i[39]),
        .I1(w_run_up_41),
        .I2(w_run_up_39),
        .O(\r_data[7]_i_1__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__39 
       (.I0(load_i[40]),
        .I1(w_run_up_42),
        .I2(w_run_up_40),
        .O(\r_data[7]_i_1__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__4 
       (.I0(load_i[5]),
        .I1(w_run_up_7),
        .I2(w_run_up_5),
        .O(\r_data[7]_i_1__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__40 
       (.I0(load_i[41]),
        .I1(w_run_up_43),
        .I2(w_run_up_41),
        .O(\r_data[7]_i_1__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__41 
       (.I0(load_i[42]),
        .I1(w_run_up_44),
        .I2(w_run_up_42),
        .O(\r_data[7]_i_1__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__42 
       (.I0(load_i[43]),
        .I1(w_run_up_45),
        .I2(w_run_up_43),
        .O(\r_data[7]_i_1__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__43 
       (.I0(load_i[44]),
        .I1(w_run_up_46),
        .I2(w_run_up_44),
        .O(\r_data[7]_i_1__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__44 
       (.I0(load_i[45]),
        .I1(w_run_up_47),
        .I2(w_run_up_45),
        .O(\r_data[7]_i_1__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__45 
       (.I0(load_i[46]),
        .I1(w_run_up_48),
        .I2(w_run_up_46),
        .O(\r_data[7]_i_1__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__46 
       (.I0(load_i[47]),
        .I1(w_run_up_49),
        .I2(w_run_up_47),
        .O(\r_data[7]_i_1__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__47 
       (.I0(load_i[48]),
        .I1(r_run_late_66),
        .I2(w_run_up_48),
        .O(\r_data[7]_i_1__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__5 
       (.I0(load_i[6]),
        .I1(w_run_up_8),
        .I2(w_run_up_6),
        .O(\r_data[7]_i_1__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__6 
       (.I0(load_i[7]),
        .I1(w_run_up_9),
        .I2(w_run_up_7),
        .O(\r_data[7]_i_1__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__7 
       (.I0(load_i[8]),
        .I1(w_run_up_10),
        .I2(w_run_up_8),
        .O(\r_data[7]_i_1__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__8 
       (.I0(load_i[9]),
        .I1(w_run_up_11),
        .I2(w_run_up_9),
        .O(\r_data[7]_i_1__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'hFE)) 
    \r_data[7]_i_1__9 
       (.I0(load_i[10]),
        .I1(w_run_up_12),
        .I2(w_run_up_10),
        .O(\r_data[7]_i_1__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair290" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2 
       (.I0(writedata_i[7]),
        .I1(readdata_o[6]),
        .I2(load_i[0]),
        .O(\r_data[7]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair286" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__0 
       (.I0(writedata_i[15]),
        .I1(readdata_o[14]),
        .I2(load_i[1]),
        .O(\r_data[7]_i_2__0_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair282" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__1 
       (.I0(writedata_i[23]),
        .I1(readdata_o[22]),
        .I2(load_i[2]),
        .O(\r_data[7]_i_2__1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair53" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__10 
       (.I0(writedata_i[95]),
        .I1(readdata_o[94]),
        .I2(load_i[11]),
        .O(\r_data[7]_i_2__10_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair57" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__11 
       (.I0(writedata_i[103]),
        .I1(readdata_o[102]),
        .I2(load_i[12]),
        .O(\r_data[7]_i_2__11_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair61" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__12 
       (.I0(writedata_i[111]),
        .I1(readdata_o[110]),
        .I2(load_i[13]),
        .O(\r_data[7]_i_2__12_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair65" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__13 
       (.I0(writedata_i[119]),
        .I1(readdata_o[118]),
        .I2(load_i[14]),
        .O(\r_data[7]_i_2__13_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair70" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__14 
       (.I0(writedata_i[127]),
        .I1(readdata_o[126]),
        .I2(load_i[15]),
        .O(\r_data[7]_i_2__14_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair74" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__15 
       (.I0(writedata_i[135]),
        .I1(readdata_o[134]),
        .I2(load_i[16]),
        .O(\r_data[7]_i_2__15_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair78" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__16 
       (.I0(writedata_i[143]),
        .I1(readdata_o[142]),
        .I2(load_i[17]),
        .O(\r_data[7]_i_2__16_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair126" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__17 
       (.I0(writedata_i[151]),
        .I1(readdata_o[150]),
        .I2(load_i[18]),
        .O(\r_data[7]_i_2__17_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair142" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__18 
       (.I0(writedata_i[159]),
        .I1(readdata_o[158]),
        .I2(load_i[19]),
        .O(\r_data[7]_i_2__18_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair90" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__19 
       (.I0(writedata_i[167]),
        .I1(readdata_o[166]),
        .I2(load_i[20]),
        .O(\r_data[7]_i_2__19_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair278" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__2 
       (.I0(writedata_i[31]),
        .I1(readdata_o[30]),
        .I2(load_i[3]),
        .O(\r_data[7]_i_2__2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair94" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__20 
       (.I0(writedata_i[175]),
        .I1(readdata_o[174]),
        .I2(load_i[21]),
        .O(\r_data[7]_i_2__20_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair99" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__21 
       (.I0(writedata_i[183]),
        .I1(readdata_o[182]),
        .I2(load_i[22]),
        .O(\r_data[7]_i_2__21_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair103" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__22 
       (.I0(writedata_i[191]),
        .I1(readdata_o[190]),
        .I2(load_i[23]),
        .O(\r_data[7]_i_2__22_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair107" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__23 
       (.I0(writedata_i[199]),
        .I1(readdata_o[198]),
        .I2(load_i[24]),
        .O(\r_data[7]_i_2__23_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair111" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__24 
       (.I0(writedata_i[207]),
        .I1(readdata_o[206]),
        .I2(load_i[25]),
        .O(\r_data[7]_i_2__24_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair115" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__25 
       (.I0(writedata_i[215]),
        .I1(readdata_o[214]),
        .I2(load_i[26]),
        .O(\r_data[7]_i_2__25_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair119" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__26 
       (.I0(writedata_i[223]),
        .I1(readdata_o[222]),
        .I2(load_i[27]),
        .O(\r_data[7]_i_2__26_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair125" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__27 
       (.I0(writedata_i[231]),
        .I1(readdata_o[230]),
        .I2(load_i[28]),
        .O(\r_data[7]_i_2__27_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair226" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__28 
       (.I0(writedata_i[239]),
        .I1(readdata_o[238]),
        .I2(load_i[29]),
        .O(\r_data[7]_i_2__28_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair232" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__29 
       (.I0(writedata_i[247]),
        .I1(readdata_o[246]),
        .I2(load_i[30]),
        .O(\r_data[7]_i_2__29_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair274" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__3 
       (.I0(writedata_i[39]),
        .I1(readdata_o[38]),
        .I2(load_i[4]),
        .O(\r_data[7]_i_2__3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair141" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__30 
       (.I0(writedata_i[255]),
        .I1(readdata_o[254]),
        .I2(load_i[31]),
        .O(\r_data[7]_i_2__30_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair246" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__31 
       (.I0(writedata_i[263]),
        .I1(readdata_o[262]),
        .I2(load_i[32]),
        .O(\r_data[7]_i_2__31_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair252" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__32 
       (.I0(writedata_i[271]),
        .I1(readdata_o[270]),
        .I2(load_i[33]),
        .O(\r_data[7]_i_2__32_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair156" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__33 
       (.I0(writedata_i[279]),
        .I1(readdata_o[278]),
        .I2(load_i[34]),
        .O(\r_data[7]_i_2__33_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair160" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__34 
       (.I0(writedata_i[287]),
        .I1(readdata_o[286]),
        .I2(load_i[35]),
        .O(\r_data[7]_i_2__34_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair164" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__35 
       (.I0(writedata_i[295]),
        .I1(readdata_o[294]),
        .I2(load_i[36]),
        .O(\r_data[7]_i_2__35_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair168" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__36 
       (.I0(writedata_i[303]),
        .I1(readdata_o[302]),
        .I2(load_i[37]),
        .O(\r_data[7]_i_2__36_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair172" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__37 
       (.I0(writedata_i[311]),
        .I1(readdata_o[310]),
        .I2(load_i[38]),
        .O(\r_data[7]_i_2__37_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair176" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__38 
       (.I0(writedata_i[319]),
        .I1(readdata_o[318]),
        .I2(load_i[39]),
        .O(\r_data[7]_i_2__38_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair180" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__39 
       (.I0(writedata_i[327]),
        .I1(readdata_o[326]),
        .I2(load_i[40]),
        .O(\r_data[7]_i_2__39_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair263" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__4 
       (.I0(writedata_i[47]),
        .I1(readdata_o[46]),
        .I2(load_i[5]),
        .O(\r_data[7]_i_2__4_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair184" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__40 
       (.I0(writedata_i[335]),
        .I1(readdata_o[334]),
        .I2(load_i[41]),
        .O(\r_data[7]_i_2__40_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair188" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__41 
       (.I0(writedata_i[343]),
        .I1(readdata_o[342]),
        .I2(load_i[42]),
        .O(\r_data[7]_i_2__41_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair192" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__42 
       (.I0(writedata_i[351]),
        .I1(readdata_o[350]),
        .I2(load_i[43]),
        .O(\r_data[7]_i_2__42_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair196" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__43 
       (.I0(writedata_i[359]),
        .I1(readdata_o[358]),
        .I2(load_i[44]),
        .O(\r_data[7]_i_2__43_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair200" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__44 
       (.I0(writedata_i[367]),
        .I1(readdata_o[366]),
        .I2(load_i[45]),
        .O(\r_data[7]_i_2__44_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair204" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__45 
       (.I0(writedata_i[375]),
        .I1(readdata_o[374]),
        .I2(load_i[46]),
        .O(\r_data[7]_i_2__45_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair208" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__46 
       (.I0(writedata_i[383]),
        .I1(readdata_o[382]),
        .I2(load_i[47]),
        .O(\r_data[7]_i_2__46_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair212" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__47 
       (.I0(writedata_i[391]),
        .I1(readdata_o[390]),
        .I2(load_i[48]),
        .O(\r_data[7]_i_2__47_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair146" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__5 
       (.I0(writedata_i[55]),
        .I1(readdata_o[54]),
        .I2(load_i[6]),
        .O(\r_data[7]_i_2__5_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair131" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__6 
       (.I0(writedata_i[63]),
        .I1(readdata_o[62]),
        .I2(load_i[7]),
        .O(\r_data[7]_i_2__6_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair88" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__7 
       (.I0(writedata_i[71]),
        .I1(readdata_o[70]),
        .I2(load_i[8]),
        .O(\r_data[7]_i_2__7_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair84" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__8 
       (.I0(writedata_i[79]),
        .I1(readdata_o[78]),
        .I2(load_i[9]),
        .O(\r_data[7]_i_2__8_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair80" *) 
  LUT3 #(
    .INIT(8'hAC)) 
    \r_data[7]_i_2__9 
       (.I0(writedata_i[87]),
        .I1(readdata_o[86]),
        .I2(load_i[10]),
        .O(\r_data[7]_i_2__9_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT3 #(
    .INIT(8'h04)) 
    r_done_i_1
       (.I0(w_run_up_49),
        .I1(\interrupt_module/r_run_delay ),
        .I2(\interrupt_module/r_swap_delay ),
        .O(r_done_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair47" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1
       (.I0(\STAGEN[1].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_1),
        .I2(readdata_o[15]),
        .I3(w_run_up_1),
        .O(r_freeze_compare_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair46" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__0
       (.I0(\STAGEN[2].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_2),
        .I2(readdata_o[23]),
        .I3(w_run_up_2),
        .O(r_freeze_compare_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair41" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__1
       (.I0(\STAGEN[3].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_3),
        .I2(readdata_o[31]),
        .I3(w_run_up_3),
        .O(r_freeze_compare_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair37" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__10
       (.I0(\STAGEN[12].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_12),
        .I2(readdata_o[103]),
        .I3(w_run_up_12),
        .O(r_freeze_compare_i_1__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair36" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__11
       (.I0(\STAGEN[13].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_13),
        .I2(readdata_o[111]),
        .I3(w_run_up_13),
        .O(r_freeze_compare_i_1__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair35" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__12
       (.I0(\STAGEN[14].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_14),
        .I2(readdata_o[119]),
        .I3(w_run_up_14),
        .O(r_freeze_compare_i_1__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair34" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__13
       (.I0(\STAGEN[15].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_15),
        .I2(readdata_o[127]),
        .I3(w_run_up_15),
        .O(r_freeze_compare_i_1__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair33" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__14
       (.I0(\STAGEN[16].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_16),
        .I2(readdata_o[135]),
        .I3(w_run_up_16),
        .O(r_freeze_compare_i_1__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair32" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__15
       (.I0(\STAGEN[17].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_17),
        .I2(readdata_o[143]),
        .I3(w_run_up_17),
        .O(r_freeze_compare_i_1__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair27" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__16
       (.I0(\STAGEN[18].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_18),
        .I2(readdata_o[151]),
        .I3(w_run_up_18),
        .O(r_freeze_compare_i_1__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair7" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__17
       (.I0(\STAGEN[19].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_19),
        .I2(readdata_o[159]),
        .I3(w_run_up_19),
        .O(r_freeze_compare_i_1__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair2" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__18
       (.I0(\STAGEN[20].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_20),
        .I2(readdata_o[167]),
        .I3(w_run_up_20),
        .O(r_freeze_compare_i_1__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair3" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__19
       (.I0(\STAGEN[21].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_21),
        .I2(readdata_o[175]),
        .I3(w_run_up_21),
        .O(r_freeze_compare_i_1__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair45" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__2
       (.I0(\STAGEN[4].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_4),
        .I2(readdata_o[39]),
        .I3(w_run_up_4),
        .O(r_freeze_compare_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair0" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__20
       (.I0(\STAGEN[22].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_22),
        .I2(readdata_o[183]),
        .I3(w_run_up_22),
        .O(r_freeze_compare_i_1__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair26" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__21
       (.I0(\STAGEN[23].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_23),
        .I2(readdata_o[191]),
        .I3(w_run_up_23),
        .O(r_freeze_compare_i_1__21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair25" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__22
       (.I0(\STAGEN[24].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_24),
        .I2(readdata_o[199]),
        .I3(w_run_up_24),
        .O(r_freeze_compare_i_1__22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair24" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__23
       (.I0(\STAGEN[25].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_25),
        .I2(readdata_o[207]),
        .I3(w_run_up_25),
        .O(r_freeze_compare_i_1__23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair23" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__24
       (.I0(\STAGEN[26].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_26),
        .I2(readdata_o[215]),
        .I3(w_run_up_26),
        .O(r_freeze_compare_i_1__24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair22" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__25
       (.I0(\STAGEN[27].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_27),
        .I2(readdata_o[223]),
        .I3(w_run_up_27),
        .O(r_freeze_compare_i_1__25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair21" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__26
       (.I0(\STAGEN[28].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_28),
        .I2(readdata_o[231]),
        .I3(w_run_up_28),
        .O(r_freeze_compare_i_1__26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair20" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__27
       (.I0(\STAGEN[29].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_29),
        .I2(readdata_o[239]),
        .I3(w_run_up_29),
        .O(r_freeze_compare_i_1__27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair19" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__28
       (.I0(\STAGEN[30].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_30),
        .I2(readdata_o[247]),
        .I3(w_run_up_30),
        .O(r_freeze_compare_i_1__28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair18" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__29
       (.I0(\STAGEN[31].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_31),
        .I2(readdata_o[255]),
        .I3(w_run_up_31),
        .O(r_freeze_compare_i_1__29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair44" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__3
       (.I0(\STAGEN[5].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_5),
        .I2(readdata_o[47]),
        .I3(w_run_up_5),
        .O(r_freeze_compare_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair17" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__30
       (.I0(\STAGEN[32].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_32),
        .I2(readdata_o[263]),
        .I3(w_run_up_32),
        .O(r_freeze_compare_i_1__30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair16" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__31
       (.I0(\STAGEN[33].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_33),
        .I2(readdata_o[271]),
        .I3(w_run_up_33),
        .O(r_freeze_compare_i_1__31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair15" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__32
       (.I0(\STAGEN[34].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_34),
        .I2(readdata_o[279]),
        .I3(w_run_up_34),
        .O(r_freeze_compare_i_1__32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair14" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__33
       (.I0(\STAGEN[35].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_35),
        .I2(readdata_o[287]),
        .I3(w_run_up_35),
        .O(r_freeze_compare_i_1__33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair13" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__34
       (.I0(\STAGEN[36].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_36),
        .I2(readdata_o[295]),
        .I3(w_run_up_36),
        .O(r_freeze_compare_i_1__34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair12" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__35
       (.I0(\STAGEN[37].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_37),
        .I2(readdata_o[303]),
        .I3(w_run_up_37),
        .O(r_freeze_compare_i_1__35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair11" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__36
       (.I0(\STAGEN[38].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_38),
        .I2(readdata_o[311]),
        .I3(w_run_up_38),
        .O(r_freeze_compare_i_1__36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair10" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__37
       (.I0(\STAGEN[39].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_39),
        .I2(readdata_o[319]),
        .I3(w_run_up_39),
        .O(r_freeze_compare_i_1__37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair9" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__38
       (.I0(\STAGEN[40].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_40),
        .I2(readdata_o[327]),
        .I3(w_run_up_40),
        .O(r_freeze_compare_i_1__38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair8" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__39
       (.I0(\STAGEN[41].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_41),
        .I2(readdata_o[335]),
        .I3(w_run_up_41),
        .O(r_freeze_compare_i_1__39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair43" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__4
       (.I0(\STAGEN[6].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_6),
        .I2(readdata_o[55]),
        .I3(w_run_up_6),
        .O(r_freeze_compare_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair1" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__40
       (.I0(\STAGEN[42].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_42),
        .I2(readdata_o[343]),
        .I3(w_run_up_42),
        .O(r_freeze_compare_i_1__40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair48" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__41
       (.I0(\STAGEN[43].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_43),
        .I2(readdata_o[351]),
        .I3(w_run_up_43),
        .O(r_freeze_compare_i_1__41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair42" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__42
       (.I0(\STAGEN[44].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_44),
        .I2(readdata_o[359]),
        .I3(w_run_up_44),
        .O(r_freeze_compare_i_1__42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair31" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__43
       (.I0(\STAGEN[45].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_45),
        .I2(readdata_o[367]),
        .I3(w_run_up_45),
        .O(r_freeze_compare_i_1__43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair30" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__44
       (.I0(\STAGEN[46].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_46),
        .I2(readdata_o[375]),
        .I3(w_run_up_46),
        .O(r_freeze_compare_i_1__44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair6" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__45
       (.I0(\STAGEN[47].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_47),
        .I2(readdata_o[383]),
        .I3(w_run_up_47),
        .O(r_freeze_compare_i_1__45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair5" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__46
       (.I0(\STAGEN[48].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_48),
        .I2(readdata_o[391]),
        .I3(w_run_up_48),
        .O(r_freeze_compare_i_1__46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair40" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__5
       (.I0(\STAGEN[7].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_7),
        .I2(readdata_o[63]),
        .I3(w_run_up_7),
        .O(r_freeze_compare_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair29" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__6
       (.I0(\STAGEN[8].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_8),
        .I2(readdata_o[71]),
        .I3(w_run_up_8),
        .O(r_freeze_compare_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair28" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__7
       (.I0(\STAGEN[9].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_9),
        .I2(readdata_o[79]),
        .I3(w_run_up_9),
        .O(r_freeze_compare_i_1__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair39" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__8
       (.I0(\STAGEN[10].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_10),
        .I2(readdata_o[87]),
        .I3(w_run_up_10),
        .O(r_freeze_compare_i_1__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair38" *) 
  LUT4 #(
    .INIT(16'hBE00)) 
    r_freeze_compare_i_1__9
       (.I0(\STAGEN[11].stage/split_module/r_freeze_compare_reg_n_0 ),
        .I1(w_bit_up_11),
        .I2(readdata_o[95]),
        .I3(w_run_up_11),
        .O(r_freeze_compare_i_1__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT4 #(
    .INIT(16'hFFF4)) 
    r_job_done_i_1
       (.I0(start_i),
        .I1(\run_module/r_job_done ),
        .I2(done_o),
        .I3(rst),
        .O(r_job_done_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1
       (.I0(\STAGEN[1].stage/split_module/r_bit1 ),
        .I1(\STAGEN[1].stage/split_module/r_compare_result ),
        .I2(\STAGEN[1].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__0
       (.I0(\STAGEN[2].stage/split_module/r_bit1 ),
        .I1(\STAGEN[2].stage/split_module/r_compare_result ),
        .I2(\STAGEN[2].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__1
       (.I0(\STAGEN[3].stage/split_module/r_bit1 ),
        .I1(\STAGEN[3].stage/split_module/r_compare_result ),
        .I2(\STAGEN[3].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__10
       (.I0(\STAGEN[12].stage/split_module/r_bit1 ),
        .I1(\STAGEN[12].stage/split_module/r_compare_result ),
        .I2(\STAGEN[12].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__11
       (.I0(\STAGEN[13].stage/split_module/r_bit1 ),
        .I1(\STAGEN[13].stage/split_module/r_compare_result ),
        .I2(\STAGEN[13].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__12
       (.I0(\STAGEN[14].stage/split_module/r_bit1 ),
        .I1(\STAGEN[14].stage/split_module/r_compare_result ),
        .I2(\STAGEN[14].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__13
       (.I0(\STAGEN[15].stage/split_module/r_bit1 ),
        .I1(\STAGEN[15].stage/split_module/r_compare_result ),
        .I2(\STAGEN[15].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__14
       (.I0(\STAGEN[16].stage/split_module/r_bit1 ),
        .I1(\STAGEN[16].stage/split_module/r_compare_result ),
        .I2(\STAGEN[16].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__15
       (.I0(\STAGEN[17].stage/split_module/r_bit1 ),
        .I1(\STAGEN[17].stage/split_module/r_compare_result ),
        .I2(\STAGEN[17].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__16
       (.I0(\STAGEN[18].stage/split_module/r_bit1 ),
        .I1(\STAGEN[18].stage/split_module/r_compare_result ),
        .I2(\STAGEN[18].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__17
       (.I0(\STAGEN[19].stage/split_module/r_bit1 ),
        .I1(\STAGEN[19].stage/split_module/r_compare_result ),
        .I2(\STAGEN[19].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__18
       (.I0(\STAGEN[20].stage/split_module/r_bit1 ),
        .I1(\STAGEN[20].stage/split_module/r_compare_result ),
        .I2(\STAGEN[20].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__19
       (.I0(\STAGEN[21].stage/split_module/r_bit1 ),
        .I1(\STAGEN[21].stage/split_module/r_compare_result ),
        .I2(\STAGEN[21].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__2
       (.I0(\STAGEN[4].stage/split_module/r_bit1 ),
        .I1(\STAGEN[4].stage/split_module/r_compare_result ),
        .I2(\STAGEN[4].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__20
       (.I0(\STAGEN[22].stage/split_module/r_bit1 ),
        .I1(\STAGEN[22].stage/split_module/r_compare_result ),
        .I2(\STAGEN[22].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__21
       (.I0(\STAGEN[23].stage/split_module/r_bit1 ),
        .I1(\STAGEN[23].stage/split_module/r_compare_result ),
        .I2(\STAGEN[23].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__22
       (.I0(\STAGEN[24].stage/split_module/r_bit1 ),
        .I1(\STAGEN[24].stage/split_module/r_compare_result ),
        .I2(\STAGEN[24].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__23
       (.I0(\STAGEN[25].stage/split_module/r_bit1 ),
        .I1(\STAGEN[25].stage/split_module/r_compare_result ),
        .I2(\STAGEN[25].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__24
       (.I0(\STAGEN[26].stage/split_module/r_bit1 ),
        .I1(\STAGEN[26].stage/split_module/r_compare_result ),
        .I2(\STAGEN[26].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__25
       (.I0(\STAGEN[27].stage/split_module/r_bit1 ),
        .I1(\STAGEN[27].stage/split_module/r_compare_result ),
        .I2(\STAGEN[27].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__26
       (.I0(\STAGEN[28].stage/split_module/r_bit1 ),
        .I1(\STAGEN[28].stage/split_module/r_compare_result ),
        .I2(\STAGEN[28].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__27
       (.I0(\STAGEN[29].stage/split_module/r_bit1 ),
        .I1(\STAGEN[29].stage/split_module/r_compare_result ),
        .I2(\STAGEN[29].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__28
       (.I0(\STAGEN[30].stage/split_module/r_bit1 ),
        .I1(\STAGEN[30].stage/split_module/r_compare_result ),
        .I2(\STAGEN[30].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__29
       (.I0(\STAGEN[31].stage/split_module/r_bit1 ),
        .I1(\STAGEN[31].stage/split_module/r_compare_result ),
        .I2(\STAGEN[31].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__3
       (.I0(\STAGEN[5].stage/split_module/r_bit1 ),
        .I1(\STAGEN[5].stage/split_module/r_compare_result ),
        .I2(\STAGEN[5].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__30
       (.I0(\STAGEN[32].stage/split_module/r_bit1 ),
        .I1(\STAGEN[32].stage/split_module/r_compare_result ),
        .I2(\STAGEN[32].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__31
       (.I0(\STAGEN[33].stage/split_module/r_bit1 ),
        .I1(\STAGEN[33].stage/split_module/r_compare_result ),
        .I2(\STAGEN[33].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__32
       (.I0(\STAGEN[34].stage/split_module/r_bit1 ),
        .I1(\STAGEN[34].stage/split_module/r_compare_result ),
        .I2(\STAGEN[34].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__33
       (.I0(\STAGEN[35].stage/split_module/r_bit1 ),
        .I1(\STAGEN[35].stage/split_module/r_compare_result ),
        .I2(\STAGEN[35].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__34
       (.I0(\STAGEN[36].stage/split_module/r_bit1 ),
        .I1(\STAGEN[36].stage/split_module/r_compare_result ),
        .I2(\STAGEN[36].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__35
       (.I0(\STAGEN[37].stage/split_module/r_bit1 ),
        .I1(\STAGEN[37].stage/split_module/r_compare_result ),
        .I2(\STAGEN[37].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__36
       (.I0(\STAGEN[38].stage/split_module/r_bit1 ),
        .I1(\STAGEN[38].stage/split_module/r_compare_result ),
        .I2(\STAGEN[38].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__37
       (.I0(\STAGEN[39].stage/split_module/r_bit1 ),
        .I1(\STAGEN[39].stage/split_module/r_compare_result ),
        .I2(\STAGEN[39].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__38
       (.I0(\STAGEN[40].stage/split_module/r_bit1 ),
        .I1(\STAGEN[40].stage/split_module/r_compare_result ),
        .I2(\STAGEN[40].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__39
       (.I0(\STAGEN[41].stage/split_module/r_bit1 ),
        .I1(\STAGEN[41].stage/split_module/r_compare_result ),
        .I2(\STAGEN[41].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__4
       (.I0(\STAGEN[6].stage/split_module/r_bit1 ),
        .I1(\STAGEN[6].stage/split_module/r_compare_result ),
        .I2(\STAGEN[6].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__40
       (.I0(\STAGEN[42].stage/split_module/r_bit1 ),
        .I1(\STAGEN[42].stage/split_module/r_compare_result ),
        .I2(\STAGEN[42].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__41
       (.I0(\STAGEN[43].stage/split_module/r_bit1 ),
        .I1(\STAGEN[43].stage/split_module/r_compare_result ),
        .I2(\STAGEN[43].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__42
       (.I0(\STAGEN[44].stage/split_module/r_bit1 ),
        .I1(\STAGEN[44].stage/split_module/r_compare_result ),
        .I2(\STAGEN[44].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__43
       (.I0(\STAGEN[45].stage/split_module/r_bit1 ),
        .I1(\STAGEN[45].stage/split_module/r_compare_result ),
        .I2(\STAGEN[45].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__44
       (.I0(\STAGEN[46].stage/split_module/r_bit1 ),
        .I1(\STAGEN[46].stage/split_module/r_compare_result ),
        .I2(\STAGEN[46].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__45
       (.I0(\STAGEN[47].stage/split_module/r_bit1 ),
        .I1(\STAGEN[47].stage/split_module/r_compare_result ),
        .I2(\STAGEN[47].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__5
       (.I0(\STAGEN[7].stage/split_module/r_bit1 ),
        .I1(\STAGEN[7].stage/split_module/r_compare_result ),
        .I2(\STAGEN[7].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__6
       (.I0(\STAGEN[8].stage/split_module/r_bit1 ),
        .I1(\STAGEN[8].stage/split_module/r_compare_result ),
        .I2(\STAGEN[8].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__7
       (.I0(\STAGEN[9].stage/split_module/r_bit1 ),
        .I1(\STAGEN[9].stage/split_module/r_compare_result ),
        .I2(\STAGEN[9].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__8
       (.I0(\STAGEN[10].stage/split_module/r_bit1 ),
        .I1(\STAGEN[10].stage/split_module/r_compare_result ),
        .I2(\STAGEN[10].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_large_bit_i_1__9
       (.I0(\STAGEN[11].stage/split_module/r_bit1 ),
        .I1(\STAGEN[11].stage/split_module/r_compare_result ),
        .I2(\STAGEN[11].stage/split_module/r_bit2 ),
        .O(r_large_bit_i_1__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT1 #(
    .INIT(2'h1)) 
    \r_pulses[0]_i_1 
       (.I0(\interrupt_module/r_pulses_reg_n_0_ ),
        .O(r_pulses0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h9)) 
    \r_pulses[1]_i_1 
       (.I0(\interrupt_module/r_pulses_reg_n_0_ ),
        .I1(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .O(r_pulses));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT3 #(
    .INIT(8'hE1)) 
    \r_pulses[2]_i_1 
       (.I0(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .I1(\interrupt_module/r_pulses_reg_n_0_ ),
        .I2(\interrupt_module/r_pulses_reg_n_0_[2] ),
        .O(\r_pulses[2]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair49" *) 
  LUT4 #(
    .INIT(16'hFE01)) 
    \r_pulses[3]_i_1 
       (.I0(\interrupt_module/r_pulses_reg_n_0_[2] ),
        .I1(\interrupt_module/r_pulses_reg_n_0_ ),
        .I2(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .I3(\interrupt_module/r_pulses_reg_n_0_[3] ),
        .O(\r_pulses[3]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair4" *) 
  LUT5 #(
    .INIT(32'hFFFE0001)) 
    \r_pulses[4]_i_1 
       (.I0(\interrupt_module/r_pulses_reg_n_0_[3] ),
        .I1(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .I2(\interrupt_module/r_pulses_reg_n_0_ ),
        .I3(\interrupt_module/r_pulses_reg_n_0_[2] ),
        .I4(\interrupt_module/r_pulses_reg_n_0_[4] ),
        .O(\r_pulses[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'hEEEEFEEE)) 
    \r_pulses[5]_i_1 
       (.I0(interrupt_o),
        .I1(rst),
        .I2(\interrupt_module/r_swap_delay ),
        .I3(\interrupt_module/r_run_delay ),
        .I4(w_run_up_49),
        .O(\r_pulses[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'h2)) 
    \r_pulses[5]_i_2 
       (.I0(\interrupt_module/r_run_delay ),
        .I1(w_run_up_49),
        .O(\r_pulses[5]_i_2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT6 #(
    .INIT(64'h00000001FFFFFFFE))
    \r_pulses[5]_i_3 
       (.I0(\interrupt_module/r_pulses_reg_n_0_[4] ),
        .I1(\interrupt_module/r_pulses_reg_n_0_[2] ),
        .I2(\interrupt_module/r_pulses_reg_n_0_ ),
        .I3(\interrupt_module/r_pulses_reg_n_0_[1] ),
        .I4(\interrupt_module/r_pulses_reg_n_0_[3] ),
        .I5(interrupt_o),
        .O(\r_pulses[5]_i_3_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_run_late_66_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run_up_49),
        .Q(r_run_late_66__0),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_run_late_66_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_run_late_66__0),
        .Q(r_run_late_66),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair213" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1
       (.I0(\STAGEN[1].stage/split_module/r_bit2 ),
        .I1(\STAGEN[1].stage/split_module/r_compare_result ),
        .I2(\STAGEN[1].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair214" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__0
       (.I0(\STAGEN[2].stage/split_module/r_bit2 ),
        .I1(\STAGEN[2].stage/split_module/r_compare_result ),
        .I2(\STAGEN[2].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__0_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair215" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__1
       (.I0(\STAGEN[3].stage/split_module/r_bit2 ),
        .I1(\STAGEN[3].stage/split_module/r_compare_result ),
        .I2(\STAGEN[3].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__1_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair227" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__10
       (.I0(\STAGEN[12].stage/split_module/r_bit2 ),
        .I1(\STAGEN[12].stage/split_module/r_compare_result ),
        .I2(\STAGEN[12].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__10_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair228" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__11
       (.I0(\STAGEN[13].stage/split_module/r_bit2 ),
        .I1(\STAGEN[13].stage/split_module/r_compare_result ),
        .I2(\STAGEN[13].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__11_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair229" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__12
       (.I0(\STAGEN[14].stage/split_module/r_bit2 ),
        .I1(\STAGEN[14].stage/split_module/r_compare_result ),
        .I2(\STAGEN[14].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__12_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair230" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__13
       (.I0(\STAGEN[15].stage/split_module/r_bit2 ),
        .I1(\STAGEN[15].stage/split_module/r_compare_result ),
        .I2(\STAGEN[15].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__13_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair231" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__14
       (.I0(\STAGEN[16].stage/split_module/r_bit2 ),
        .I1(\STAGEN[16].stage/split_module/r_compare_result ),
        .I2(\STAGEN[16].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__14_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair233" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__15
       (.I0(\STAGEN[17].stage/split_module/r_bit2 ),
        .I1(\STAGEN[17].stage/split_module/r_compare_result ),
        .I2(\STAGEN[17].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__15_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair234" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__16
       (.I0(\STAGEN[18].stage/split_module/r_bit2 ),
        .I1(\STAGEN[18].stage/split_module/r_compare_result ),
        .I2(\STAGEN[18].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__16_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair235" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__17
       (.I0(\STAGEN[19].stage/split_module/r_bit2 ),
        .I1(\STAGEN[19].stage/split_module/r_compare_result ),
        .I2(\STAGEN[19].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__17_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair236" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__18
       (.I0(\STAGEN[20].stage/split_module/r_bit2 ),
        .I1(\STAGEN[20].stage/split_module/r_compare_result ),
        .I2(\STAGEN[20].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__18_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair237" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__19
       (.I0(\STAGEN[21].stage/split_module/r_bit2 ),
        .I1(\STAGEN[21].stage/split_module/r_compare_result ),
        .I2(\STAGEN[21].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__19_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair216" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__2
       (.I0(\STAGEN[4].stage/split_module/r_bit2 ),
        .I1(\STAGEN[4].stage/split_module/r_compare_result ),
        .I2(\STAGEN[4].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__2_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair239" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__20
       (.I0(\STAGEN[22].stage/split_module/r_bit2 ),
        .I1(\STAGEN[22].stage/split_module/r_compare_result ),
        .I2(\STAGEN[22].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__20_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair240" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__21
       (.I0(\STAGEN[23].stage/split_module/r_bit2 ),
        .I1(\STAGEN[23].stage/split_module/r_compare_result ),
        .I2(\STAGEN[23].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__21_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair241" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__22
       (.I0(\STAGEN[24].stage/split_module/r_bit2 ),
        .I1(\STAGEN[24].stage/split_module/r_compare_result ),
        .I2(\STAGEN[24].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__22_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair242" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__23
       (.I0(\STAGEN[25].stage/split_module/r_bit2 ),
        .I1(\STAGEN[25].stage/split_module/r_compare_result ),
        .I2(\STAGEN[25].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__23_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair244" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__24
       (.I0(\STAGEN[26].stage/split_module/r_bit2 ),
        .I1(\STAGEN[26].stage/split_module/r_compare_result ),
        .I2(\STAGEN[26].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__24_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair245" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__25
       (.I0(\STAGEN[27].stage/split_module/r_bit2 ),
        .I1(\STAGEN[27].stage/split_module/r_compare_result ),
        .I2(\STAGEN[27].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__25_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair247" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__26
       (.I0(\STAGEN[28].stage/split_module/r_bit2 ),
        .I1(\STAGEN[28].stage/split_module/r_compare_result ),
        .I2(\STAGEN[28].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__26_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair248" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__27
       (.I0(\STAGEN[29].stage/split_module/r_bit2 ),
        .I1(\STAGEN[29].stage/split_module/r_compare_result ),
        .I2(\STAGEN[29].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__27_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair249" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__28
       (.I0(\STAGEN[30].stage/split_module/r_bit2 ),
        .I1(\STAGEN[30].stage/split_module/r_compare_result ),
        .I2(\STAGEN[30].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__28_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair250" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__29
       (.I0(\STAGEN[31].stage/split_module/r_bit2 ),
        .I1(\STAGEN[31].stage/split_module/r_compare_result ),
        .I2(\STAGEN[31].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__29_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair217" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__3
       (.I0(\STAGEN[5].stage/split_module/r_bit2 ),
        .I1(\STAGEN[5].stage/split_module/r_compare_result ),
        .I2(\STAGEN[5].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__3_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair251" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__30
       (.I0(\STAGEN[32].stage/split_module/r_bit2 ),
        .I1(\STAGEN[32].stage/split_module/r_compare_result ),
        .I2(\STAGEN[32].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__30_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair253" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__31
       (.I0(\STAGEN[33].stage/split_module/r_bit2 ),
        .I1(\STAGEN[33].stage/split_module/r_compare_result ),
        .I2(\STAGEN[33].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__31_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair254" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__32
       (.I0(\STAGEN[34].stage/split_module/r_bit2 ),
        .I1(\STAGEN[34].stage/split_module/r_compare_result ),
        .I2(\STAGEN[34].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__32_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair255" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__33
       (.I0(\STAGEN[35].stage/split_module/r_bit2 ),
        .I1(\STAGEN[35].stage/split_module/r_compare_result ),
        .I2(\STAGEN[35].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__33_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair256" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__34
       (.I0(\STAGEN[36].stage/split_module/r_bit2 ),
        .I1(\STAGEN[36].stage/split_module/r_compare_result ),
        .I2(\STAGEN[36].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__34_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair257" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__35
       (.I0(\STAGEN[37].stage/split_module/r_bit2 ),
        .I1(\STAGEN[37].stage/split_module/r_compare_result ),
        .I2(\STAGEN[37].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__35_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair259" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__36
       (.I0(\STAGEN[38].stage/split_module/r_bit2 ),
        .I1(\STAGEN[38].stage/split_module/r_compare_result ),
        .I2(\STAGEN[38].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__36_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair260" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__37
       (.I0(\STAGEN[39].stage/split_module/r_bit2 ),
        .I1(\STAGEN[39].stage/split_module/r_compare_result ),
        .I2(\STAGEN[39].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__37_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair261" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__38
       (.I0(\STAGEN[40].stage/split_module/r_bit2 ),
        .I1(\STAGEN[40].stage/split_module/r_compare_result ),
        .I2(\STAGEN[40].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__38_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair262" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__39
       (.I0(\STAGEN[41].stage/split_module/r_bit2 ),
        .I1(\STAGEN[41].stage/split_module/r_compare_result ),
        .I2(\STAGEN[41].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__39_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair219" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__4
       (.I0(\STAGEN[6].stage/split_module/r_bit2 ),
        .I1(\STAGEN[6].stage/split_module/r_compare_result ),
        .I2(\STAGEN[6].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__4_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair264" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__40
       (.I0(\STAGEN[42].stage/split_module/r_bit2 ),
        .I1(\STAGEN[42].stage/split_module/r_compare_result ),
        .I2(\STAGEN[42].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__40_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair265" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__41
       (.I0(\STAGEN[43].stage/split_module/r_bit2 ),
        .I1(\STAGEN[43].stage/split_module/r_compare_result ),
        .I2(\STAGEN[43].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__41_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair267" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__42
       (.I0(\STAGEN[44].stage/split_module/r_bit2 ),
        .I1(\STAGEN[44].stage/split_module/r_compare_result ),
        .I2(\STAGEN[44].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__42_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair269" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__43
       (.I0(\STAGEN[45].stage/split_module/r_bit2 ),
        .I1(\STAGEN[45].stage/split_module/r_compare_result ),
        .I2(\STAGEN[45].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__43_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair271" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__44
       (.I0(\STAGEN[46].stage/split_module/r_bit2 ),
        .I1(\STAGEN[46].stage/split_module/r_compare_result ),
        .I2(\STAGEN[46].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__44_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair272" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__45
       (.I0(\STAGEN[47].stage/split_module/r_bit2 ),
        .I1(\STAGEN[47].stage/split_module/r_compare_result ),
        .I2(\STAGEN[47].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__45_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__46
       (.I0(\STAGEN[48].stage/split_module/r_bit2 ),
        .I1(\STAGEN[48].stage/split_module/r_compare_result ),
        .I2(\STAGEN[48].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__46_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair220" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__5
       (.I0(\STAGEN[7].stage/split_module/r_bit2 ),
        .I1(\STAGEN[7].stage/split_module/r_compare_result ),
        .I2(\STAGEN[7].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__5_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair221" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__6
       (.I0(\STAGEN[8].stage/split_module/r_bit2 ),
        .I1(\STAGEN[8].stage/split_module/r_compare_result ),
        .I2(\STAGEN[8].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__6_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair222" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__7
       (.I0(\STAGEN[9].stage/split_module/r_bit2 ),
        .I1(\STAGEN[9].stage/split_module/r_compare_result ),
        .I2(\STAGEN[9].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__7_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair224" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__8
       (.I0(\STAGEN[10].stage/split_module/r_bit2 ),
        .I1(\STAGEN[10].stage/split_module/r_compare_result ),
        .I2(\STAGEN[10].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__8_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair225" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    r_small_bit_i_1__9
       (.I0(\STAGEN[11].stage/split_module/r_bit2 ),
        .I1(\STAGEN[11].stage/split_module/r_compare_result ),
        .I2(\STAGEN[11].stage/split_module/r_bit1 ),
        .O(r_small_bit_i_1__9_n_0));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1 
       (.I0(\STAGEN[2].stage/split_module/p_0_in ),
        .I1(\STAGEN[2].stage/split_module/r_compare_result ),
        .O(\STAGEN[2].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__0 
       (.I0(\STAGEN[3].stage/split_module/p_0_in ),
        .I1(\STAGEN[3].stage/split_module/r_compare_result ),
        .O(\STAGEN[3].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__1 
       (.I0(\STAGEN[4].stage/split_module/p_0_in ),
        .I1(\STAGEN[4].stage/split_module/r_compare_result ),
        .O(\STAGEN[4].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__10 
       (.I0(\STAGEN[13].stage/split_module/p_0_in ),
        .I1(\STAGEN[13].stage/split_module/r_compare_result ),
        .O(\STAGEN[13].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__11 
       (.I0(\STAGEN[14].stage/split_module/p_0_in ),
        .I1(\STAGEN[14].stage/split_module/r_compare_result ),
        .O(\STAGEN[14].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__12 
       (.I0(\STAGEN[15].stage/split_module/p_0_in ),
        .I1(\STAGEN[15].stage/split_module/r_compare_result ),
        .O(\STAGEN[15].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__13 
       (.I0(\STAGEN[16].stage/split_module/p_0_in ),
        .I1(\STAGEN[16].stage/split_module/r_compare_result ),
        .O(\STAGEN[16].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__14 
       (.I0(\STAGEN[17].stage/split_module/p_0_in ),
        .I1(\STAGEN[17].stage/split_module/r_compare_result ),
        .O(\STAGEN[17].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__15 
       (.I0(\STAGEN[18].stage/split_module/p_0_in ),
        .I1(\STAGEN[18].stage/split_module/r_compare_result ),
        .O(\STAGEN[18].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__16 
       (.I0(\STAGEN[19].stage/split_module/p_0_in ),
        .I1(\STAGEN[19].stage/split_module/r_compare_result ),
        .O(\STAGEN[19].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__17 
       (.I0(\STAGEN[20].stage/split_module/p_0_in ),
        .I1(\STAGEN[20].stage/split_module/r_compare_result ),
        .O(\STAGEN[20].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__18 
       (.I0(\STAGEN[21].stage/split_module/p_0_in ),
        .I1(\STAGEN[21].stage/split_module/r_compare_result ),
        .O(\STAGEN[21].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__19 
       (.I0(\STAGEN[22].stage/split_module/p_0_in ),
        .I1(\STAGEN[22].stage/split_module/r_compare_result ),
        .O(\STAGEN[22].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__2 
       (.I0(\STAGEN[5].stage/split_module/p_0_in ),
        .I1(\STAGEN[5].stage/split_module/r_compare_result ),
        .O(\STAGEN[5].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__20 
       (.I0(\STAGEN[23].stage/split_module/p_0_in ),
        .I1(\STAGEN[23].stage/split_module/r_compare_result ),
        .O(\STAGEN[23].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__21 
       (.I0(\STAGEN[24].stage/split_module/p_0_in ),
        .I1(\STAGEN[24].stage/split_module/r_compare_result ),
        .O(\STAGEN[24].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__22 
       (.I0(\STAGEN[25].stage/split_module/p_0_in ),
        .I1(\STAGEN[25].stage/split_module/r_compare_result ),
        .O(\STAGEN[25].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__23 
       (.I0(\STAGEN[26].stage/split_module/p_0_in ),
        .I1(\STAGEN[26].stage/split_module/r_compare_result ),
        .O(\STAGEN[26].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__24 
       (.I0(\STAGEN[27].stage/split_module/p_0_in ),
        .I1(\STAGEN[27].stage/split_module/r_compare_result ),
        .O(\STAGEN[27].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__25 
       (.I0(\STAGEN[28].stage/split_module/p_0_in ),
        .I1(\STAGEN[28].stage/split_module/r_compare_result ),
        .O(\STAGEN[28].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__26 
       (.I0(\STAGEN[29].stage/split_module/p_0_in ),
        .I1(\STAGEN[29].stage/split_module/r_compare_result ),
        .O(\STAGEN[29].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__27 
       (.I0(\STAGEN[30].stage/split_module/p_0_in ),
        .I1(\STAGEN[30].stage/split_module/r_compare_result ),
        .O(\STAGEN[30].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__28 
       (.I0(\STAGEN[31].stage/split_module/p_0_in ),
        .I1(\STAGEN[31].stage/split_module/r_compare_result ),
        .O(\STAGEN[31].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__29 
       (.I0(\STAGEN[32].stage/split_module/p_0_in ),
        .I1(\STAGEN[32].stage/split_module/r_compare_result ),
        .O(\STAGEN[32].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__3 
       (.I0(\STAGEN[6].stage/split_module/p_0_in ),
        .I1(\STAGEN[6].stage/split_module/r_compare_result ),
        .O(\STAGEN[6].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__30 
       (.I0(\STAGEN[33].stage/split_module/p_0_in ),
        .I1(\STAGEN[33].stage/split_module/r_compare_result ),
        .O(\STAGEN[33].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__31 
       (.I0(\STAGEN[34].stage/split_module/p_0_in ),
        .I1(\STAGEN[34].stage/split_module/r_compare_result ),
        .O(\STAGEN[34].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__32 
       (.I0(\STAGEN[35].stage/split_module/p_0_in ),
        .I1(\STAGEN[35].stage/split_module/r_compare_result ),
        .O(\STAGEN[35].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__33 
       (.I0(\STAGEN[36].stage/split_module/p_0_in ),
        .I1(\STAGEN[36].stage/split_module/r_compare_result ),
        .O(\STAGEN[36].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__34 
       (.I0(\STAGEN[37].stage/split_module/p_0_in ),
        .I1(\STAGEN[37].stage/split_module/r_compare_result ),
        .O(\STAGEN[37].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__35 
       (.I0(\STAGEN[38].stage/split_module/p_0_in ),
        .I1(\STAGEN[38].stage/split_module/r_compare_result ),
        .O(\STAGEN[38].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__36 
       (.I0(\STAGEN[39].stage/split_module/p_0_in ),
        .I1(\STAGEN[39].stage/split_module/r_compare_result ),
        .O(\STAGEN[39].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__37 
       (.I0(\STAGEN[40].stage/split_module/p_0_in ),
        .I1(\STAGEN[40].stage/split_module/r_compare_result ),
        .O(\STAGEN[40].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__38 
       (.I0(\STAGEN[41].stage/split_module/p_0_in ),
        .I1(\STAGEN[41].stage/split_module/r_compare_result ),
        .O(\STAGEN[41].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__39 
       (.I0(\STAGEN[42].stage/split_module/p_0_in ),
        .I1(\STAGEN[42].stage/split_module/r_compare_result ),
        .O(\STAGEN[42].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__4 
       (.I0(\STAGEN[7].stage/split_module/p_0_in ),
        .I1(\STAGEN[7].stage/split_module/r_compare_result ),
        .O(\STAGEN[7].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__40 
       (.I0(\STAGEN[43].stage/split_module/p_0_in ),
        .I1(\STAGEN[43].stage/split_module/r_compare_result ),
        .O(\STAGEN[43].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__41 
       (.I0(\STAGEN[44].stage/split_module/p_0_in ),
        .I1(\STAGEN[44].stage/split_module/r_compare_result ),
        .O(\STAGEN[44].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__42 
       (.I0(\STAGEN[45].stage/split_module/p_0_in ),
        .I1(\STAGEN[45].stage/split_module/r_compare_result ),
        .O(\STAGEN[45].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__43 
       (.I0(\STAGEN[46].stage/split_module/p_0_in ),
        .I1(\STAGEN[46].stage/split_module/r_compare_result ),
        .O(\STAGEN[46].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__44 
       (.I0(\STAGEN[47].stage/split_module/p_0_in ),
        .I1(\STAGEN[47].stage/split_module/r_compare_result ),
        .O(\STAGEN[47].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__45 
       (.I0(\STAGEN[48].stage/split_module/p_0_in ),
        .I1(\STAGEN[48].stage/split_module/r_compare_result ),
        .O(\STAGEN[48].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__5 
       (.I0(\STAGEN[8].stage/split_module/p_0_in ),
        .I1(\STAGEN[8].stage/split_module/r_compare_result ),
        .O(\STAGEN[8].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__6 
       (.I0(\STAGEN[9].stage/split_module/p_0_in ),
        .I1(\STAGEN[9].stage/split_module/r_compare_result ),
        .O(\STAGEN[9].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__7 
       (.I0(\STAGEN[10].stage/split_module/p_0_in ),
        .I1(\STAGEN[10].stage/split_module/r_compare_result ),
        .O(\STAGEN[10].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__8 
       (.I0(\STAGEN[11].stage/split_module/p_0_in ),
        .I1(\STAGEN[11].stage/split_module/r_compare_result ),
        .O(\STAGEN[11].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \r_swap[1]_i_1__9 
       (.I0(\STAGEN[12].stage/split_module/p_0_in ),
        .I1(\STAGEN[12].stage/split_module/r_compare_result ),
        .O(\STAGEN[12].stage/split_module/p_1_out ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* srl_bus_name = "bubblesort_0/\r_value_66_reg " *) 
  (* srl_name = "bubblesort_0/\r_value_66_reg[0]_srl2 " *) 
  SRL16E #(
    .INIT(16'h0000),
    .IS_CLK_INVERTED(1'b0)) 
    \r_value_66_reg[0]_srl2 
       (.A0(\<const1>__0__0 ),
        .A1(\<const0>__0__0 ),
        .A2(\<const0>__0__0 ),
        .A3(\<const0>__0__0 ),
        .CE(\<const1>__0__0 ),
        .CLK(clk),
        .D(r_value_66_reg),
        .Q(\r_value_66_reg[0]_srl2_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair273" *) 
  LUT3 #(
    .INIT(8'hB8)) 
    \r_value_66_reg[0]_srl2_i_1 
       (.I0(\STAGEN[48].stage/split_module/r_bit1 ),
        .I1(\STAGEN[48].stage/split_module/r_compare_result ),
        .I2(\STAGEN[48].stage/split_module/r_bit2 ),
        .O(r_value_66_reg));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \r_value_66_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\r_value_66_reg[0]_srl2_n_0 ),
        .Q(r_value_66),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  LUT5 #(
    .INIT(32'h00002022)) 
    \run_module/r_count[0]_i_1 
       (.I0(p_2_in[0]),
        .I1(rst),
        .I2(w_run),
        .I3(\run_module/r_job_done ),
        .I4(start_i),
        .O(\run_module/r_count ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[10]_i_1 
       (.I0(p_2_in[10]),
        .I1(start_i),
        .O(\run_module/r_count[10]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[11]_i_1 
       (.I0(p_2_in[11]),
        .I1(start_i),
        .O(\run_module/r_count[11]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair294" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[4]_i_1 
       (.I0(p_2_in[4]),
        .I1(start_i),
        .O(\run_module/r_count[4]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair295" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[5]_i_1 
       (.I0(p_2_in[5]),
        .I1(start_i),
        .O(\run_module/r_count[5]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[6]_i_1 
       (.I0(p_2_in[6]),
        .I1(start_i),
        .O(\run_module/r_count[6]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[7]_i_1 
       (.I0(p_2_in[7]),
        .I1(start_i),
        .O(\run_module/r_count[7]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair297" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[8]_i_1 
       (.I0(p_2_in[8]),
        .I1(start_i),
        .O(\run_module/r_count[8]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* SOFT_HLUTNM = "soft_lutpair296" *) 
  LUT2 #(
    .INIT(4'hE)) 
    \run_module/r_count[9]_i_1 
       (.I0(p_2_in[9]),
        .I1(start_i),
        .O(\run_module/r_count[9]_i_1_n_0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[0] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count ),
        .Q(w_run),
        .R(\<const0>__0__0 ));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[10] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[10]_i_1_n_0 ),
        .Q(p_2_in[11]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[11] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[11]_i_1_n_0 ),
        .Q(p_2_in[0]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[1] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(w_run),
        .Q(p_2_in[2]),
        .R(r_count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[2] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_2_in[2]),
        .Q(p_2_in[3]),
        .R(r_count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[3] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(p_2_in[3]),
        .Q(p_2_in[4]),
        .R(r_count));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[4] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[4]_i_1_n_0 ),
        .Q(p_2_in[5]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[5] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[5]_i_1_n_0 ),
        .Q(p_2_in[6]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[6] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[6]_i_1_n_0 ),
        .Q(p_2_in[7]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[7] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[7]_i_1_n_0 ),
        .Q(p_2_in[8]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[8] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[8]_i_1_n_0 ),
        .Q(p_2_in[9]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_count_reg[9] 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(\run_module/r_count[9]_i_1_n_0 ),
        .Q(p_2_in[10]),
        .R(rst));
  (* BOX_TYPE = "PRIMITIVE" *) 
  (* STRUCTURAL_NETLIST = "yes" *) 
  FDRE #(
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .IS_R_INVERTED(1'b0)) 
    \run_module/r_job_done_reg 
       (.C(clk),
        .CE(\<const1>__0__0 ),
        .D(r_job_done_i_1_n_0),
        .Q(\run_module/r_job_done ),
        .R(\<const0>__0__0 ));
endmodule
